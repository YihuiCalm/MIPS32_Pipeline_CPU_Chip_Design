// Created by ihdl
module MIPS32_CPU_top ( clk, rst_n, instruction, inst_address );
  input [31:0] instruction;
  output [31:0] inst_address;
  input clk, rst_n;
  wire   inst_ID2EX_reg_N170, inst_ID2EX_reg_N169, inst_ID2EX_reg_N168,
         inst_ID2EX_reg_N167, inst_ID2EX_reg_N166, inst_ID2EX_reg_N139,
         inst_ID2EX_reg_N138, inst_ID2EX_reg_N137, inst_ID2EX_reg_N136,
         inst_ID2EX_reg_N135, inst_ID2EX_reg_N134, inst_ID2EX_reg_N117,
         inst_ID2EX_reg_N116, inst_ID2EX_reg_N115, inst_ID2EX_reg_N114,
         inst_ID2EX_reg_N113, inst_ID2EX_reg_N112, inst_ID2EX_reg_N111,
         inst_ID2EX_reg_N110, inst_ID2EX_reg_N109, inst_ID2EX_reg_N108,
         inst_ID2EX_reg_N107, inst_ID2EX_reg_N106, inst_ID2EX_reg_N105,
         inst_ID2EX_reg_N104, inst_ID2EX_reg_N103, inst_ID2EX_reg_N102,
         inst_ID2EX_reg_N101, inst_ID2EX_reg_N100, inst_ID2EX_reg_N99,
         inst_ID2EX_reg_N98, inst_ID2EX_reg_N97, inst_ID2EX_reg_N96,
         inst_ID2EX_reg_N95, inst_ID2EX_reg_N94, inst_ID2EX_reg_N93,
         inst_ID2EX_reg_N92, inst_ID2EX_reg_N91, inst_ID2EX_reg_N90,
         inst_ID2EX_reg_N89, inst_ID2EX_reg_N88, inst_ID2EX_reg_N87,
         inst_ID2EX_reg_N86, inst_ID2EX_reg_N85, inst_ID2EX_reg_N84,
         inst_ID2EX_reg_N83, inst_ID2EX_reg_N82, inst_ID2EX_reg_N81,
         inst_ID2EX_reg_N80, inst_ID2EX_reg_N79, inst_ID2EX_reg_N78,
         inst_ID2EX_reg_N77, inst_ID2EX_reg_N76, inst_ID2EX_reg_N75,
         inst_ID2EX_reg_N74, inst_ID2EX_reg_N73, inst_ID2EX_reg_N72,
         inst_ID2EX_reg_N71, inst_ID2EX_reg_N70, inst_ID2EX_reg_N69,
         inst_ID2EX_reg_N68, inst_ID2EX_reg_N67, inst_ID2EX_reg_N66,
         inst_ID2EX_reg_N65, inst_ID2EX_reg_N64, inst_ID2EX_reg_N63,
         inst_ID2EX_reg_N62, inst_ID2EX_reg_N61, inst_ID2EX_reg_N60,
         inst_ID2EX_reg_N59, inst_ID2EX_reg_N58, inst_ID2EX_reg_N57,
         inst_ID2EX_reg_N56, inst_ID2EX_reg_N55, inst_ID2EX_reg_N54,
         inst_ID2EX_reg_N53, inst_ID2EX_reg_N52, inst_ID2EX_reg_N51,
         inst_ID2EX_reg_N50, inst_ID2EX_reg_N49, inst_ID2EX_reg_N48,
         inst_ID2EX_reg_N47, inst_ID2EX_reg_N46, inst_ID2EX_reg_N45,
         inst_ID2EX_reg_N44, inst_ID2EX_reg_N43, inst_ID2EX_reg_N42,
         inst_ID2EX_reg_N41, inst_ID2EX_reg_N40, inst_ID2EX_reg_N39,
         inst_ID2EX_reg_N38, inst_ID2EX_reg_N37, inst_ID2EX_reg_N36,
         inst_ID2EX_reg_N35, inst_ID2EX_reg_N34, inst_ID2EX_reg_N33,
         inst_ID2EX_reg_N32, inst_ID2EX_reg_N31, inst_ID2EX_reg_N30,
         inst_ID2EX_reg_N29, inst_ID2EX_reg_N28, inst_ID2EX_reg_N27,
         inst_ID2EX_reg_N26, inst_ID2EX_reg_N25, inst_ID2EX_reg_N24,
         inst_ID2EX_reg_N23, inst_ID2EX_reg_N22, inst_ID2EX_reg_N21,
         inst_ID2EX_reg_N20, inst_ID2EX_reg_N19, inst_ID2EX_reg_N18,
         inst_ID2EX_reg_N17, inst_ID2EX_reg_N16, inst_ID2EX_reg_N15,
         inst_ID2EX_reg_N14, inst_ID2EX_reg_N13, inst_ID2EX_reg_N12,
         inst_ID2EX_reg_N11, inst_ID2EX_reg_N10, inst_ID2EX_reg_N9,
         inst_ID2EX_reg_N8, inst_ID2EX_reg_N7, inst_ID2EX_reg_N6,
         inst_ID2EX_reg_N5, inst_ID2EX_reg_N4, inst_ID2EX_reg_N3,
         inst_EX2MEM_reg_N133, inst_EX2MEM_reg_N132, inst_EX2MEM_reg_N131,
         inst_EX2MEM_reg_N130, inst_EX2MEM_reg_N129, inst_EX2MEM_reg_N128,
         inst_EX2MEM_reg_N127, inst_EX2MEM_reg_N126, inst_EX2MEM_reg_N125,
         inst_EX2MEM_reg_N124, inst_EX2MEM_reg_N123, inst_EX2MEM_reg_N122,
         inst_EX2MEM_reg_N121, inst_EX2MEM_reg_N120, inst_EX2MEM_reg_N119,
         inst_EX2MEM_reg_N118, inst_EX2MEM_reg_N117, inst_EX2MEM_reg_N116,
         inst_EX2MEM_reg_N115, inst_EX2MEM_reg_N114, inst_EX2MEM_reg_N113,
         inst_EX2MEM_reg_N112, inst_EX2MEM_reg_N111, inst_EX2MEM_reg_N110,
         inst_EX2MEM_reg_N109, inst_EX2MEM_reg_N108, inst_EX2MEM_reg_N107,
         inst_EX2MEM_reg_N106, inst_EX2MEM_reg_N105, inst_EX2MEM_reg_N104,
         inst_EX2MEM_reg_N103, inst_EX2MEM_reg_N102, inst_EX2MEM_reg_N101,
         inst_EX2MEM_reg_N100, inst_EX2MEM_reg_N99, inst_EX2MEM_reg_N98,
         inst_EX2MEM_reg_N97, inst_EX2MEM_reg_N96, inst_EX2MEM_reg_N95,
         inst_EX2MEM_reg_N94, inst_EX2MEM_reg_N93, inst_EX2MEM_reg_N92,
         inst_EX2MEM_reg_N91, inst_EX2MEM_reg_N90, inst_EX2MEM_reg_N89,
         inst_EX2MEM_reg_N88, inst_EX2MEM_reg_N87, inst_EX2MEM_reg_N86,
         inst_EX2MEM_reg_N85, inst_EX2MEM_reg_N84, inst_EX2MEM_reg_N83,
         inst_EX2MEM_reg_N82, inst_EX2MEM_reg_N81, inst_EX2MEM_reg_N80,
         inst_EX2MEM_reg_N79, inst_EX2MEM_reg_N78, inst_EX2MEM_reg_N77,
         inst_EX2MEM_reg_N76, inst_EX2MEM_reg_N75, inst_EX2MEM_reg_N74,
         inst_EX2MEM_reg_N73, inst_EX2MEM_reg_N72, inst_EX2MEM_reg_N71,
         inst_EX2MEM_reg_N70, inst_EX2MEM_reg_N69, inst_EX2MEM_reg_N68,
         inst_EX2MEM_reg_N67, inst_EX2MEM_reg_N66, inst_EX2MEM_reg_N65,
         inst_EX2MEM_reg_N64, inst_EX2MEM_reg_N63, inst_EX2MEM_reg_N62,
         inst_EX2MEM_reg_N61, inst_EX2MEM_reg_N60, inst_EX2MEM_reg_N59,
         inst_EX2MEM_reg_N58, inst_EX2MEM_reg_N57, inst_EX2MEM_reg_N56,
         inst_EX2MEM_reg_N55, inst_EX2MEM_reg_N54, inst_EX2MEM_reg_N53,
         inst_EX2MEM_reg_N52, inst_EX2MEM_reg_N51, inst_EX2MEM_reg_N50,
         inst_EX2MEM_reg_N49, inst_EX2MEM_reg_N48, inst_EX2MEM_reg_N47,
         inst_EX2MEM_reg_N46, inst_EX2MEM_reg_N45, inst_EX2MEM_reg_N44,
         inst_EX2MEM_reg_N43, inst_EX2MEM_reg_N42, inst_EX2MEM_reg_N41,
         inst_EX2MEM_reg_N40, inst_EX2MEM_reg_N39, inst_EX2MEM_reg_N38,
         inst_EX2MEM_reg_N37, inst_EX2MEM_reg_N36, inst_EX2MEM_reg_N35,
         inst_EX2MEM_reg_N34, inst_EX2MEM_reg_N33, inst_EX2MEM_reg_N32,
         inst_EX2MEM_reg_N31, inst_EX2MEM_reg_N30, inst_EX2MEM_reg_N29,
         inst_EX2MEM_reg_N28, inst_EX2MEM_reg_N27, inst_EX2MEM_reg_N26,
         inst_EX2MEM_reg_N25, inst_EX2MEM_reg_N24, inst_EX2MEM_reg_N23,
         inst_EX2MEM_reg_N22, inst_EX2MEM_reg_N21, inst_EX2MEM_reg_N20,
         inst_EX2MEM_reg_N19, inst_EX2MEM_reg_N18, inst_EX2MEM_reg_N17,
         inst_EX2MEM_reg_N16, inst_EX2MEM_reg_N15, inst_EX2MEM_reg_N14,
         inst_EX2MEM_reg_N13, inst_EX2MEM_reg_N12, inst_EX2MEM_reg_N11,
         inst_EX2MEM_reg_N10, inst_EX2MEM_reg_N9, inst_EX2MEM_reg_N8,
         inst_EX2MEM_reg_N7, inst_EX2MEM_reg_N6, inst_EX2MEM_reg_N5,
         inst_EX2MEM_reg_N4, inst_EX2MEM_reg_N3, u_MEM2WB_reg_N75,
         u_MEM2WB_reg_N74, u_MEM2WB_reg_N73, u_MEM2WB_reg_N72,
         u_MEM2WB_reg_N71, u_MEM2WB_reg_N70, u_MEM2WB_reg_N69,
         u_MEM2WB_reg_N68, u_MEM2WB_reg_N67, u_MEM2WB_reg_N66,
         u_MEM2WB_reg_N65, u_MEM2WB_reg_N64, u_MEM2WB_reg_N63,
         u_MEM2WB_reg_N62, u_MEM2WB_reg_N61, u_MEM2WB_reg_N60,
         u_MEM2WB_reg_N59, u_MEM2WB_reg_N58, u_MEM2WB_reg_N57,
         u_MEM2WB_reg_N56, u_MEM2WB_reg_N55, u_MEM2WB_reg_N54,
         u_MEM2WB_reg_N53, u_MEM2WB_reg_N52, u_MEM2WB_reg_N51,
         u_MEM2WB_reg_N50, u_MEM2WB_reg_N49, u_MEM2WB_reg_N48,
         u_MEM2WB_reg_N47, u_MEM2WB_reg_N46, u_MEM2WB_reg_N45,
         u_MEM2WB_reg_N44, u_MEM2WB_reg_N43, u_MEM2WB_reg_N42,
         u_MEM2WB_reg_N41, u_MEM2WB_reg_N40, u_MEM2WB_reg_N39,
         u_MEM2WB_reg_N38, u_MEM2WB_reg_N37, u_MEM2WB_reg_N36,
         u_MEM2WB_reg_N35, u_MEM2WB_reg_N34, u_MEM2WB_reg_N33,
         u_MEM2WB_reg_N32, u_MEM2WB_reg_N31, u_MEM2WB_reg_N30,
         u_MEM2WB_reg_N29, u_MEM2WB_reg_N28, u_MEM2WB_reg_N27,
         u_MEM2WB_reg_N26, u_MEM2WB_reg_N25, u_MEM2WB_reg_N24,
         u_MEM2WB_reg_N23, u_MEM2WB_reg_N22, u_MEM2WB_reg_N21,
         u_MEM2WB_reg_N20, u_MEM2WB_reg_N19, u_MEM2WB_reg_N18,
         u_MEM2WB_reg_N17, u_MEM2WB_reg_N16, u_MEM2WB_reg_N15,
         u_MEM2WB_reg_N14, u_MEM2WB_reg_N13, u_MEM2WB_reg_N12,
         u_MEM2WB_reg_N11, u_MEM2WB_reg_N10, u_MEM2WB_reg_N9, u_MEM2WB_reg_N8,
         u_MEM2WB_reg_N7, u_MEM2WB_reg_N6, u_MEM2WB_reg_N5, u_MEM2WB_reg_N4,
         u_MEM2WB_reg_N3, n2183, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528;
  wire   [31:0] instruction_ID;
  wire   [31:0] inst_addr_ID;
  wire   [4:0] reg_write_address_WB;
  wire   [3:0] op_type_EX;
  wire   [31:2] inst_addr_EX;
  wire   [31:0] reg_read_data_1_EX;
  wire   [31:0] reg_read_data_2_EX;
  wire   [15:0] jump_inst_addr_EX;
  wire   [4:0] read_register_1_EX;
  wire   [4:0] read_register_2_EX;
  wire   [4:0] reg_write_address_MEM;
  wire   [31:0] alu_result_MEM;
  wire   [1:0] shifted_address_EX;
  wire   [3:0] op_type_MEM;
  wire   [31:0] shifted_address_MEM;
  wire   [31:0] write_mem_data_MEM;
  wire   [25:0] jump_inst_addr_MEM;
  wire   [3:0] op_type_WB;
  wire   [31:0] mem_read_data_WB;
  wire   [31:0] alu_result_WB;
  wire   [255:0] inst_register_registers;
  wire   [255:0] inst_data_MEM_data;

  DFFPOSX1 inst_data_MEM_data_reg_7__31_ ( .D(n2726), .CLK(clk), .Q(
        inst_data_MEM_data[255]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_31_ ( .D(u_MEM2WB_reg_N38), .CLK(clk), 
        .Q(mem_read_data_WB[31]) );
  DFFPOSX1 inst_register_registers_reg_0__31_ ( .D(n2246), .CLK(clk), .Q(
        inst_register_registers[31]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_31_ ( .D(inst_ID2EX_reg_N70), .CLK(
        clk), .Q(reg_read_data_1_EX[31]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_31_ ( .D(inst_EX2MEM_reg_N70), .CLK(
        clk), .Q(alu_result_MEM[31]) );
  DFFPOSX1 inst_ID2EX_reg_op_type_reg_3_ ( .D(inst_ID2EX_reg_N6), .CLK(clk), 
        .Q(op_type_EX[3]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_31_ ( .D(n2790), .CLK(clk), .Q(
        instruction_ID[31]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_30_ ( .D(n2789), .CLK(clk), .Q(
        instruction_ID[30]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_29_ ( .D(n2788), .CLK(clk), .Q(
        instruction_ID[29]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_28_ ( .D(n2787), .CLK(clk), .Q(
        instruction_ID[28]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_27_ ( .D(n2786), .CLK(clk), .Q(
        instruction_ID[27]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_26_ ( .D(n2785), .CLK(clk), .Q(
        instruction_ID[26]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_25_ ( .D(n2784), .CLK(clk), .Q(
        instruction_ID[25]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_addr_reg_4_ ( .D(inst_ID2EX_reg_N170), 
        .CLK(clk), .Q(read_register_1_EX[4]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_24_ ( .D(n2783), .CLK(clk), .Q(
        instruction_ID[24]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_addr_reg_3_ ( .D(inst_ID2EX_reg_N169), 
        .CLK(clk), .Q(read_register_1_EX[3]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_23_ ( .D(n2782), .CLK(clk), .Q(
        instruction_ID[23]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_addr_reg_2_ ( .D(inst_ID2EX_reg_N168), 
        .CLK(clk), .Q(read_register_1_EX[2]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_22_ ( .D(n2781), .CLK(clk), .Q(
        instruction_ID[22]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_addr_reg_1_ ( .D(inst_ID2EX_reg_N167), 
        .CLK(clk), .Q(read_register_1_EX[1]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_21_ ( .D(n2780), .CLK(clk), .Q(
        instruction_ID[21]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_addr_reg_0_ ( .D(inst_ID2EX_reg_N166), 
        .CLK(clk), .Q(read_register_1_EX[0]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_20_ ( .D(n2779), .CLK(clk), .Q(
        instruction_ID[20]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_addr_reg_4_ ( .D(inst_ID2EX_reg_N139), 
        .CLK(clk), .Q(read_register_2_EX[4]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_19_ ( .D(n2778), .CLK(clk), .Q(
        instruction_ID[19]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_addr_reg_3_ ( .D(inst_ID2EX_reg_N138), 
        .CLK(clk), .Q(read_register_2_EX[3]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_18_ ( .D(n2777), .CLK(clk), .Q(
        instruction_ID[18]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_addr_reg_2_ ( .D(inst_ID2EX_reg_N137), 
        .CLK(clk), .Q(read_register_2_EX[2]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_17_ ( .D(n2776), .CLK(clk), .Q(
        instruction_ID[17]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_addr_reg_1_ ( .D(inst_ID2EX_reg_N136), 
        .CLK(clk), .Q(read_register_2_EX[1]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_16_ ( .D(n2775), .CLK(clk), .Q(
        instruction_ID[16]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_addr_reg_0_ ( .D(inst_ID2EX_reg_N135), 
        .CLK(clk), .Q(read_register_2_EX[0]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_15_ ( .D(n2774), .CLK(clk), .Q(
        instruction_ID[15]) );
  DFFPOSX1 inst_ID2EX_reg_jump_address_reg_15_ ( .D(inst_ID2EX_reg_N134), 
        .CLK(clk), .Q(jump_inst_addr_EX[15]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_14_ ( .D(n2773), .CLK(clk), .Q(
        instruction_ID[14]) );
  DFFPOSX1 inst_ID2EX_reg_jump_address_reg_14_ ( .D(inst_ID2EX_reg_N117), 
        .CLK(clk), .Q(jump_inst_addr_EX[14]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_13_ ( .D(n2772), .CLK(clk), .Q(
        instruction_ID[13]) );
  DFFPOSX1 inst_ID2EX_reg_jump_address_reg_13_ ( .D(inst_ID2EX_reg_N116), 
        .CLK(clk), .Q(jump_inst_addr_EX[13]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_12_ ( .D(n2771), .CLK(clk), .Q(
        instruction_ID[12]) );
  DFFPOSX1 inst_ID2EX_reg_jump_address_reg_12_ ( .D(inst_ID2EX_reg_N115), 
        .CLK(clk), .Q(jump_inst_addr_EX[12]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_11_ ( .D(n2770), .CLK(clk), .Q(
        instruction_ID[11]) );
  DFFPOSX1 inst_ID2EX_reg_jump_address_reg_11_ ( .D(inst_ID2EX_reg_N114), 
        .CLK(clk), .Q(jump_inst_addr_EX[11]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_10_ ( .D(n2769), .CLK(clk), .Q(
        instruction_ID[10]) );
  DFFPOSX1 inst_ID2EX_reg_jump_address_reg_10_ ( .D(inst_ID2EX_reg_N113), 
        .CLK(clk), .Q(jump_inst_addr_EX[10]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_9_ ( .D(n2768), .CLK(clk), .Q(
        instruction_ID[9]) );
  DFFPOSX1 inst_ID2EX_reg_jump_address_reg_9_ ( .D(inst_ID2EX_reg_N112), .CLK(
        clk), .Q(jump_inst_addr_EX[9]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_8_ ( .D(n2767), .CLK(clk), .Q(
        instruction_ID[8]) );
  DFFPOSX1 inst_ID2EX_reg_jump_address_reg_8_ ( .D(inst_ID2EX_reg_N111), .CLK(
        clk), .Q(jump_inst_addr_EX[8]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_7_ ( .D(n2766), .CLK(clk), .Q(
        instruction_ID[7]) );
  DFFPOSX1 inst_ID2EX_reg_jump_address_reg_7_ ( .D(inst_ID2EX_reg_N110), .CLK(
        clk), .Q(jump_inst_addr_EX[7]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_6_ ( .D(n2765), .CLK(clk), .Q(
        instruction_ID[6]) );
  DFFPOSX1 inst_ID2EX_reg_jump_address_reg_6_ ( .D(inst_ID2EX_reg_N109), .CLK(
        clk), .Q(jump_inst_addr_EX[6]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_5_ ( .D(n2764), .CLK(clk), .Q(
        instruction_ID[5]) );
  DFFPOSX1 inst_ID2EX_reg_jump_address_reg_5_ ( .D(inst_ID2EX_reg_N108), .CLK(
        clk), .Q(jump_inst_addr_EX[5]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_4_ ( .D(n2763), .CLK(clk), .Q(
        instruction_ID[4]) );
  DFFPOSX1 inst_ID2EX_reg_jump_address_reg_4_ ( .D(inst_ID2EX_reg_N107), .CLK(
        clk), .Q(jump_inst_addr_EX[4]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_3_ ( .D(n2762), .CLK(clk), .Q(
        instruction_ID[3]) );
  DFFPOSX1 inst_ID2EX_reg_jump_address_reg_3_ ( .D(inst_ID2EX_reg_N106), .CLK(
        clk), .Q(jump_inst_addr_EX[3]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_2_ ( .D(n2761), .CLK(clk), .Q(
        instruction_ID[2]) );
  DFFPOSX1 inst_ID2EX_reg_jump_address_reg_2_ ( .D(inst_ID2EX_reg_N105), .CLK(
        clk), .Q(jump_inst_addr_EX[2]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_1_ ( .D(n2760), .CLK(clk), .Q(
        instruction_ID[1]) );
  DFFPOSX1 inst_ID2EX_reg_jump_address_reg_1_ ( .D(inst_ID2EX_reg_N104), .CLK(
        clk), .Q(jump_inst_addr_EX[1]) );
  DFFPOSX1 inst_IF2ID_reg_instruction_reg_0_ ( .D(n2759), .CLK(clk), .Q(
        instruction_ID[0]) );
  DFFPOSX1 inst_ID2EX_reg_jump_address_reg_0_ ( .D(inst_ID2EX_reg_N103), .CLK(
        clk), .Q(jump_inst_addr_EX[0]) );
  DFFPOSX1 inst_ID2EX_reg_op_type_reg_1_ ( .D(inst_ID2EX_reg_N4), .CLK(clk), 
        .Q(op_type_EX[1]) );
  DFFPOSX1 inst_ID2EX_reg_op_type_reg_0_ ( .D(inst_ID2EX_reg_N3), .CLK(clk), 
        .Q(op_type_EX[0]) );
  DFFPOSX1 inst_ID2EX_reg_op_type_reg_2_ ( .D(inst_ID2EX_reg_N5), .CLK(clk), 
        .Q(op_type_EX[2]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_0_ ( .D(inst_EX2MEM_reg_N108), 
        .CLK(clk), .Q(jump_inst_addr_MEM[0]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_1_ ( .D(inst_EX2MEM_reg_N109), 
        .CLK(clk), .Q(jump_inst_addr_MEM[1]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_2_ ( .D(inst_EX2MEM_reg_N110), 
        .CLK(clk), .Q(jump_inst_addr_MEM[2]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_3_ ( .D(inst_EX2MEM_reg_N111), 
        .CLK(clk), .Q(jump_inst_addr_MEM[3]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_4_ ( .D(inst_EX2MEM_reg_N112), 
        .CLK(clk), .Q(jump_inst_addr_MEM[4]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_5_ ( .D(inst_EX2MEM_reg_N113), 
        .CLK(clk), .Q(jump_inst_addr_MEM[5]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_6_ ( .D(inst_EX2MEM_reg_N114), 
        .CLK(clk), .Q(jump_inst_addr_MEM[6]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_7_ ( .D(inst_EX2MEM_reg_N115), 
        .CLK(clk), .Q(jump_inst_addr_MEM[7]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_8_ ( .D(inst_EX2MEM_reg_N116), 
        .CLK(clk), .Q(jump_inst_addr_MEM[8]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_9_ ( .D(inst_EX2MEM_reg_N117), 
        .CLK(clk), .Q(jump_inst_addr_MEM[9]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_10_ ( .D(inst_EX2MEM_reg_N118), 
        .CLK(clk), .Q(jump_inst_addr_MEM[10]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_11_ ( .D(inst_EX2MEM_reg_N119), 
        .CLK(clk), .Q(jump_inst_addr_MEM[11]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_12_ ( .D(inst_EX2MEM_reg_N120), 
        .CLK(clk), .Q(jump_inst_addr_MEM[12]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_13_ ( .D(inst_EX2MEM_reg_N121), 
        .CLK(clk), .Q(jump_inst_addr_MEM[13]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_14_ ( .D(inst_EX2MEM_reg_N122), 
        .CLK(clk), .Q(jump_inst_addr_MEM[14]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_15_ ( .D(inst_EX2MEM_reg_N123), 
        .CLK(clk), .Q(jump_inst_addr_MEM[15]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_16_ ( .D(inst_EX2MEM_reg_N124), 
        .CLK(clk), .Q(jump_inst_addr_MEM[16]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_17_ ( .D(inst_EX2MEM_reg_N125), 
        .CLK(clk), .Q(jump_inst_addr_MEM[17]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_18_ ( .D(inst_EX2MEM_reg_N126), 
        .CLK(clk), .Q(jump_inst_addr_MEM[18]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_19_ ( .D(inst_EX2MEM_reg_N127), 
        .CLK(clk), .Q(jump_inst_addr_MEM[19]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_20_ ( .D(inst_EX2MEM_reg_N128), 
        .CLK(clk), .Q(jump_inst_addr_MEM[20]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_21_ ( .D(inst_EX2MEM_reg_N129), 
        .CLK(clk), .Q(jump_inst_addr_MEM[21]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_22_ ( .D(inst_EX2MEM_reg_N130), 
        .CLK(clk), .Q(jump_inst_addr_MEM[22]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_23_ ( .D(inst_EX2MEM_reg_N131), 
        .CLK(clk), .Q(jump_inst_addr_MEM[23]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_24_ ( .D(inst_EX2MEM_reg_N132), 
        .CLK(clk), .Q(jump_inst_addr_MEM[24]) );
  DFFPOSX1 inst_EX2MEM_reg_jump_address_reg_25_ ( .D(inst_EX2MEM_reg_N133), 
        .CLK(clk), .Q(jump_inst_addr_MEM[25]) );
  DFFPOSX1 inst_EX2MEM_reg_write_reg_address_reg_0_ ( .D(inst_EX2MEM_reg_N103), 
        .CLK(clk), .Q(reg_write_address_MEM[0]) );
  DFFPOSX1 inst_EX2MEM_reg_write_reg_address_reg_1_ ( .D(inst_EX2MEM_reg_N104), 
        .CLK(clk), .Q(reg_write_address_MEM[1]) );
  DFFPOSX1 inst_EX2MEM_reg_write_reg_address_reg_2_ ( .D(inst_EX2MEM_reg_N105), 
        .CLK(clk), .Q(reg_write_address_MEM[2]) );
  DFFPOSX1 inst_EX2MEM_reg_write_reg_address_reg_3_ ( .D(inst_EX2MEM_reg_N106), 
        .CLK(clk), .Q(reg_write_address_MEM[3]) );
  DFFPOSX1 inst_EX2MEM_reg_write_reg_address_reg_4_ ( .D(inst_EX2MEM_reg_N107), 
        .CLK(clk), .Q(reg_write_address_MEM[4]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_0_ ( .D(inst_EX2MEM_reg_N7), 
        .CLK(clk), .Q(shifted_address_MEM[0]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_1_ ( .D(inst_EX2MEM_reg_N8), 
        .CLK(clk), .Q(shifted_address_MEM[1]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_2_ ( .D(inst_EX2MEM_reg_N9), 
        .CLK(clk), .Q(shifted_address_MEM[2]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_3_ ( .D(inst_EX2MEM_reg_N10), 
        .CLK(clk), .Q(shifted_address_MEM[3]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_4_ ( .D(inst_EX2MEM_reg_N11), 
        .CLK(clk), .Q(shifted_address_MEM[4]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_5_ ( .D(inst_EX2MEM_reg_N12), 
        .CLK(clk), .Q(shifted_address_MEM[5]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_6_ ( .D(inst_EX2MEM_reg_N13), 
        .CLK(clk), .Q(shifted_address_MEM[6]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_7_ ( .D(inst_EX2MEM_reg_N14), 
        .CLK(clk), .Q(shifted_address_MEM[7]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_8_ ( .D(inst_EX2MEM_reg_N15), 
        .CLK(clk), .Q(shifted_address_MEM[8]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_9_ ( .D(inst_EX2MEM_reg_N16), 
        .CLK(clk), .Q(shifted_address_MEM[9]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_10_ ( .D(inst_EX2MEM_reg_N17), 
        .CLK(clk), .Q(shifted_address_MEM[10]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_11_ ( .D(inst_EX2MEM_reg_N18), 
        .CLK(clk), .Q(shifted_address_MEM[11]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_12_ ( .D(inst_EX2MEM_reg_N19), 
        .CLK(clk), .Q(shifted_address_MEM[12]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_13_ ( .D(inst_EX2MEM_reg_N20), 
        .CLK(clk), .Q(shifted_address_MEM[13]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_14_ ( .D(inst_EX2MEM_reg_N21), 
        .CLK(clk), .Q(shifted_address_MEM[14]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_15_ ( .D(inst_EX2MEM_reg_N22), 
        .CLK(clk), .Q(shifted_address_MEM[15]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_16_ ( .D(inst_EX2MEM_reg_N23), 
        .CLK(clk), .Q(shifted_address_MEM[16]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_17_ ( .D(inst_EX2MEM_reg_N24), 
        .CLK(clk), .Q(shifted_address_MEM[17]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_18_ ( .D(inst_EX2MEM_reg_N25), 
        .CLK(clk), .Q(shifted_address_MEM[18]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_19_ ( .D(inst_EX2MEM_reg_N26), 
        .CLK(clk), .Q(shifted_address_MEM[19]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_20_ ( .D(inst_EX2MEM_reg_N27), 
        .CLK(clk), .Q(shifted_address_MEM[20]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_21_ ( .D(inst_EX2MEM_reg_N28), 
        .CLK(clk), .Q(shifted_address_MEM[21]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_22_ ( .D(inst_EX2MEM_reg_N29), 
        .CLK(clk), .Q(shifted_address_MEM[22]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_23_ ( .D(inst_EX2MEM_reg_N30), 
        .CLK(clk), .Q(shifted_address_MEM[23]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_24_ ( .D(inst_EX2MEM_reg_N31), 
        .CLK(clk), .Q(shifted_address_MEM[24]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_25_ ( .D(inst_EX2MEM_reg_N32), 
        .CLK(clk), .Q(shifted_address_MEM[25]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_26_ ( .D(inst_EX2MEM_reg_N33), 
        .CLK(clk), .Q(shifted_address_MEM[26]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_27_ ( .D(inst_EX2MEM_reg_N34), 
        .CLK(clk), .Q(shifted_address_MEM[27]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_28_ ( .D(inst_EX2MEM_reg_N35), 
        .CLK(clk), .Q(shifted_address_MEM[28]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_29_ ( .D(inst_EX2MEM_reg_N36), 
        .CLK(clk), .Q(shifted_address_MEM[29]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_30_ ( .D(inst_EX2MEM_reg_N37), 
        .CLK(clk), .Q(shifted_address_MEM[30]) );
  DFFPOSX1 inst_EX2MEM_reg_shifted_address_reg_31_ ( .D(inst_EX2MEM_reg_N38), 
        .CLK(clk), .Q(shifted_address_MEM[31]) );
  DFFPOSX1 inst_EX2MEM_reg_op_type_reg_0_ ( .D(inst_EX2MEM_reg_N3), .CLK(clk), 
        .Q(op_type_MEM[0]) );
  DFFPOSX1 inst_EX2MEM_reg_op_type_reg_1_ ( .D(inst_EX2MEM_reg_N4), .CLK(clk), 
        .Q(op_type_MEM[1]) );
  DFFPOSX1 inst_EX2MEM_reg_op_type_reg_2_ ( .D(inst_EX2MEM_reg_N5), .CLK(clk), 
        .Q(op_type_MEM[2]) );
  DFFPOSX1 inst_EX2MEM_reg_op_type_reg_3_ ( .D(inst_EX2MEM_reg_N6), .CLK(clk), 
        .Q(op_type_MEM[3]) );
  DFFPOSX1 u_MEM2WB_reg_write_reg_address_reg_0_ ( .D(u_MEM2WB_reg_N71), .CLK(
        clk), .Q(reg_write_address_WB[0]) );
  DFFPOSX1 u_MEM2WB_reg_write_reg_address_reg_1_ ( .D(u_MEM2WB_reg_N72), .CLK(
        clk), .Q(reg_write_address_WB[1]) );
  DFFPOSX1 u_MEM2WB_reg_write_reg_address_reg_2_ ( .D(u_MEM2WB_reg_N73), .CLK(
        clk), .Q(reg_write_address_WB[2]) );
  DFFPOSX1 u_MEM2WB_reg_write_reg_address_reg_3_ ( .D(u_MEM2WB_reg_N74), .CLK(
        clk), .Q(reg_write_address_WB[3]) );
  DFFPOSX1 u_MEM2WB_reg_write_reg_address_reg_4_ ( .D(u_MEM2WB_reg_N75), .CLK(
        clk), .Q(reg_write_address_WB[4]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_31_ ( .D(u_MEM2WB_reg_N70), .CLK(clk), 
        .Q(alu_result_WB[31]) );
  DFFPOSX1 u_MEM2WB_reg_op_type_reg_0_ ( .D(u_MEM2WB_reg_N3), .CLK(clk), .Q(
        op_type_WB[0]) );
  DFFPOSX1 u_MEM2WB_reg_op_type_reg_1_ ( .D(u_MEM2WB_reg_N4), .CLK(clk), .Q(
        op_type_WB[1]) );
  DFFPOSX1 u_MEM2WB_reg_op_type_reg_2_ ( .D(u_MEM2WB_reg_N5), .CLK(clk), .Q(
        op_type_WB[2]) );
  DFFPOSX1 u_MEM2WB_reg_op_type_reg_3_ ( .D(u_MEM2WB_reg_N6), .CLK(clk), .Q(
        op_type_WB[3]) );
  DFFPOSX1 inst_register_registers_reg_6__31_ ( .D(n2440), .CLK(clk), .Q(
        inst_register_registers[223]) );
  DFFPOSX1 inst_register_registers_reg_7__31_ ( .D(n2314), .CLK(clk), .Q(
        inst_register_registers[255]) );
  DFFPOSX1 inst_register_registers_reg_3__31_ ( .D(n2343), .CLK(clk), .Q(
        inst_register_registers[127]) );
  DFFPOSX1 inst_register_registers_reg_2__31_ ( .D(n2310), .CLK(clk), .Q(
        inst_register_registers[95]) );
  DFFPOSX1 inst_register_registers_reg_4__31_ ( .D(n2375), .CLK(clk), .Q(
        inst_register_registers[159]) );
  DFFPOSX1 inst_register_registers_reg_5__31_ ( .D(n2407), .CLK(clk), .Q(
        inst_register_registers[191]) );
  DFFPOSX1 inst_register_registers_reg_1__31_ ( .D(n2278), .CLK(clk), .Q(
        inst_register_registers[63]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_31_ ( .D(inst_ID2EX_reg_N102), .CLK(
        clk), .Q(reg_read_data_2_EX[31]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_31_ ( .D(inst_EX2MEM_reg_N102), 
        .CLK(clk), .Q(write_mem_data_MEM[31]) );
  DFFPOSX1 inst_register_registers_reg_6__30_ ( .D(n2415), .CLK(clk), .Q(
        inst_register_registers[222]) );
  DFFPOSX1 inst_register_registers_reg_7__30_ ( .D(n2414), .CLK(clk), .Q(
        inst_register_registers[254]) );
  DFFPOSX1 inst_register_registers_reg_5__30_ ( .D(n2376), .CLK(clk), .Q(
        inst_register_registers[190]) );
  DFFPOSX1 inst_register_registers_reg_4__30_ ( .D(n2344), .CLK(clk), .Q(
        inst_register_registers[158]) );
  DFFPOSX1 inst_register_registers_reg_3__30_ ( .D(n2315), .CLK(clk), .Q(
        inst_register_registers[126]) );
  DFFPOSX1 inst_register_registers_reg_2__30_ ( .D(n2279), .CLK(clk), .Q(
        inst_register_registers[94]) );
  DFFPOSX1 inst_register_registers_reg_1__30_ ( .D(n2247), .CLK(clk), .Q(
        inst_register_registers[62]) );
  DFFPOSX1 inst_register_registers_reg_0__30_ ( .D(n2215), .CLK(clk), .Q(
        inst_register_registers[30]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_30_ ( .D(inst_ID2EX_reg_N101), .CLK(
        clk), .Q(reg_read_data_2_EX[30]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_30_ ( .D(inst_EX2MEM_reg_N101), 
        .CLK(clk), .Q(write_mem_data_MEM[30]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_30_ ( .D(inst_ID2EX_reg_N69), .CLK(
        clk), .Q(reg_read_data_1_EX[30]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_30_ ( .D(inst_EX2MEM_reg_N69), .CLK(
        clk), .Q(alu_result_MEM[30]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_30_ ( .D(u_MEM2WB_reg_N69), .CLK(clk), 
        .Q(alu_result_WB[30]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_0_ ( .D(inst_EX2MEM_reg_N39), .CLK(
        clk), .Q(alu_result_MEM[0]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_0_ ( .D(u_MEM2WB_reg_N39), .CLK(clk), 
        .Q(alu_result_WB[0]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__31_ ( .D(n2690), .CLK(clk), .Q(
        inst_data_MEM_data[63]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__30_ ( .D(n2659), .CLK(clk), .Q(
        inst_data_MEM_data[62]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_2_ ( .D(u_MEM2WB_reg_N9), .CLK(clk), .Q(
        mem_read_data_WB[2]) );
  DFFPOSX1 inst_register_registers_reg_7__2_ ( .D(n2467), .CLK(clk), .Q(
        inst_register_registers[226]) );
  DFFPOSX1 inst_register_registers_reg_6__2_ ( .D(n2410), .CLK(clk), .Q(
        inst_register_registers[194]) );
  DFFPOSX1 inst_register_registers_reg_5__2_ ( .D(n2404), .CLK(clk), .Q(
        inst_register_registers[162]) );
  DFFPOSX1 inst_register_registers_reg_4__2_ ( .D(n2372), .CLK(clk), .Q(
        inst_register_registers[130]) );
  DFFPOSX1 inst_register_registers_reg_3__2_ ( .D(n2313), .CLK(clk), .Q(
        inst_register_registers[98]) );
  DFFPOSX1 inst_register_registers_reg_2__2_ ( .D(n2307), .CLK(clk), .Q(
        inst_register_registers[66]) );
  DFFPOSX1 inst_register_registers_reg_1__2_ ( .D(n2275), .CLK(clk), .Q(
        inst_register_registers[34]) );
  DFFPOSX1 inst_register_registers_reg_0__2_ ( .D(n2243), .CLK(clk), .Q(
        inst_register_registers[2]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_2_ ( .D(inst_ID2EX_reg_N73), .CLK(clk), .Q(reg_read_data_2_EX[2]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_2_ ( .D(inst_EX2MEM_reg_N73), 
        .CLK(clk), .Q(write_mem_data_MEM[2]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__2_ ( .D(n2687), .CLK(clk), .Q(
        inst_data_MEM_data[34]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_2_ ( .D(inst_ID2EX_reg_N41), .CLK(clk), .Q(reg_read_data_1_EX[2]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_2_ ( .D(inst_EX2MEM_reg_N41), .CLK(
        clk), .Q(alu_result_MEM[2]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_2_ ( .D(u_MEM2WB_reg_N41), .CLK(clk), 
        .Q(alu_result_WB[2]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__2_ ( .D(n2725), .CLK(clk), .Q(
        inst_data_MEM_data[98]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__1_ ( .D(n2723), .CLK(clk), .Q(
        inst_data_MEM_data[97]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_1_ ( .D(u_MEM2WB_reg_N8), .CLK(clk), .Q(
        mem_read_data_WB[1]) );
  DFFPOSX1 inst_register_registers_reg_7__1_ ( .D(n2468), .CLK(clk), .Q(
        inst_register_registers[225]) );
  DFFPOSX1 inst_register_registers_reg_6__1_ ( .D(n2411), .CLK(clk), .Q(
        inst_register_registers[193]) );
  DFFPOSX1 inst_register_registers_reg_5__1_ ( .D(n2405), .CLK(clk), .Q(
        inst_register_registers[161]) );
  DFFPOSX1 inst_register_registers_reg_4__1_ ( .D(n2373), .CLK(clk), .Q(
        inst_register_registers[129]) );
  DFFPOSX1 inst_register_registers_reg_3__1_ ( .D(n2311), .CLK(clk), .Q(
        inst_register_registers[97]) );
  DFFPOSX1 inst_register_registers_reg_2__1_ ( .D(n2308), .CLK(clk), .Q(
        inst_register_registers[65]) );
  DFFPOSX1 inst_register_registers_reg_1__1_ ( .D(n2276), .CLK(clk), .Q(
        inst_register_registers[33]) );
  DFFPOSX1 inst_register_registers_reg_0__1_ ( .D(n2244), .CLK(clk), .Q(
        inst_register_registers[1]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_1_ ( .D(inst_ID2EX_reg_N72), .CLK(clk), .Q(reg_read_data_2_EX[1]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_1_ ( .D(inst_EX2MEM_reg_N72), 
        .CLK(clk), .Q(write_mem_data_MEM[1]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__1_ ( .D(n2688), .CLK(clk), .Q(
        inst_data_MEM_data[33]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_1_ ( .D(inst_ID2EX_reg_N40), .CLK(clk), .Q(reg_read_data_1_EX[1]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_1_ ( .D(inst_EX2MEM_reg_N40), .CLK(
        clk), .Q(alu_result_MEM[1]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_1_ ( .D(u_MEM2WB_reg_N40), .CLK(clk), 
        .Q(alu_result_WB[1]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__31_ ( .D(n2722), .CLK(clk), .Q(
        inst_data_MEM_data[95]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__1_ ( .D(n2720), .CLK(clk), .Q(
        inst_data_MEM_data[65]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__2_ ( .D(n2719), .CLK(clk), .Q(
        inst_data_MEM_data[66]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__30_ ( .D(n2691), .CLK(clk), .Q(
        inst_data_MEM_data[94]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__30_ ( .D(n2626), .CLK(clk), .Q(
        inst_data_MEM_data[254]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__1_ ( .D(n2524), .CLK(clk), .Q(
        inst_data_MEM_data[225]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__2_ ( .D(n2523), .CLK(clk), .Q(
        inst_data_MEM_data[226]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__1_ ( .D(n2623), .CLK(clk), .Q(
        inst_data_MEM_data[193]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__2_ ( .D(n2622), .CLK(clk), .Q(
        inst_data_MEM_data[194]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__31_ ( .D(n2496), .CLK(clk), .Q(
        inst_data_MEM_data[223]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__30_ ( .D(n2471), .CLK(clk), .Q(
        inst_data_MEM_data[222]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__31_ ( .D(n2658), .CLK(clk), .Q(
        inst_data_MEM_data[31]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__1_ ( .D(n2656), .CLK(clk), .Q(
        inst_data_MEM_data[1]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__2_ ( .D(n2655), .CLK(clk), .Q(
        inst_data_MEM_data[2]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__30_ ( .D(n2627), .CLK(clk), .Q(
        inst_data_MEM_data[30]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__31_ ( .D(n2619), .CLK(clk), .Q(
        inst_data_MEM_data[191]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__1_ ( .D(n2617), .CLK(clk), .Q(
        inst_data_MEM_data[161]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__2_ ( .D(n2616), .CLK(clk), .Q(
        inst_data_MEM_data[162]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__30_ ( .D(n2588), .CLK(clk), .Q(
        inst_data_MEM_data[190]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__31_ ( .D(n2587), .CLK(clk), .Q(
        inst_data_MEM_data[159]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__0_ ( .D(n2586), .CLK(clk), .Q(
        inst_data_MEM_data[128]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_0_ ( .D(u_MEM2WB_reg_N7), .CLK(clk), .Q(
        mem_read_data_WB[0]) );
  DFFPOSX1 inst_register_registers_reg_7__0_ ( .D(n2469), .CLK(clk), .Q(
        inst_register_registers[224]) );
  DFFPOSX1 inst_register_registers_reg_6__0_ ( .D(n2412), .CLK(clk), .Q(
        inst_register_registers[192]) );
  DFFPOSX1 inst_register_registers_reg_5__0_ ( .D(n2406), .CLK(clk), .Q(
        inst_register_registers[160]) );
  DFFPOSX1 inst_register_registers_reg_4__0_ ( .D(n2374), .CLK(clk), .Q(
        inst_register_registers[128]) );
  DFFPOSX1 inst_register_registers_reg_3__0_ ( .D(n2312), .CLK(clk), .Q(
        inst_register_registers[96]) );
  DFFPOSX1 inst_register_registers_reg_2__0_ ( .D(n2309), .CLK(clk), .Q(
        inst_register_registers[64]) );
  DFFPOSX1 inst_register_registers_reg_1__0_ ( .D(n2277), .CLK(clk), .Q(
        inst_register_registers[32]) );
  DFFPOSX1 inst_register_registers_reg_0__0_ ( .D(n2245), .CLK(clk), .Q(
        inst_register_registers[0]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_0_ ( .D(inst_ID2EX_reg_N71), .CLK(clk), .Q(reg_read_data_2_EX[0]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_0_ ( .D(inst_EX2MEM_reg_N71), 
        .CLK(clk), .Q(write_mem_data_MEM[0]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__0_ ( .D(n2721), .CLK(clk), .Q(
        inst_data_MEM_data[64]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__0_ ( .D(n2657), .CLK(clk), .Q(
        inst_data_MEM_data[0]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__0_ ( .D(n2624), .CLK(clk), .Q(
        inst_data_MEM_data[192]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__0_ ( .D(n2724), .CLK(clk), .Q(
        inst_data_MEM_data[96]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__0_ ( .D(n2689), .CLK(clk), .Q(
        inst_data_MEM_data[32]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__0_ ( .D(n2618), .CLK(clk), .Q(
        inst_data_MEM_data[160]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__0_ ( .D(n2525), .CLK(clk), .Q(
        inst_data_MEM_data[224]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_0_ ( .D(inst_ID2EX_reg_N39), .CLK(clk), .Q(reg_read_data_1_EX[0]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__1_ ( .D(n2585), .CLK(clk), .Q(
        inst_data_MEM_data[129]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__2_ ( .D(n2584), .CLK(clk), .Q(
        inst_data_MEM_data[130]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__30_ ( .D(n2556), .CLK(clk), .Q(
        inst_data_MEM_data[158]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__31_ ( .D(n2555), .CLK(clk), .Q(
        inst_data_MEM_data[127]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__30_ ( .D(n2527), .CLK(clk), .Q(
        inst_data_MEM_data[126]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_3_ ( .D(u_MEM2WB_reg_N10), .CLK(clk), 
        .Q(mem_read_data_WB[3]) );
  DFFPOSX1 inst_register_registers_reg_7__3_ ( .D(n2466), .CLK(clk), .Q(
        inst_register_registers[227]) );
  DFFPOSX1 inst_register_registers_reg_6__3_ ( .D(n2409), .CLK(clk), .Q(
        inst_register_registers[195]) );
  DFFPOSX1 inst_register_registers_reg_5__3_ ( .D(n2403), .CLK(clk), .Q(
        inst_register_registers[163]) );
  DFFPOSX1 inst_register_registers_reg_4__3_ ( .D(n2371), .CLK(clk), .Q(
        inst_register_registers[131]) );
  DFFPOSX1 inst_register_registers_reg_3__3_ ( .D(n2342), .CLK(clk), .Q(
        inst_register_registers[99]) );
  DFFPOSX1 inst_register_registers_reg_2__3_ ( .D(n2306), .CLK(clk), .Q(
        inst_register_registers[67]) );
  DFFPOSX1 inst_register_registers_reg_1__3_ ( .D(n2274), .CLK(clk), .Q(
        inst_register_registers[35]) );
  DFFPOSX1 inst_register_registers_reg_0__3_ ( .D(n2242), .CLK(clk), .Q(
        inst_register_registers[3]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_3_ ( .D(inst_ID2EX_reg_N74), .CLK(clk), .Q(reg_read_data_2_EX[3]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_3_ ( .D(inst_EX2MEM_reg_N74), 
        .CLK(clk), .Q(write_mem_data_MEM[3]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__3_ ( .D(n2718), .CLK(clk), .Q(
        inst_data_MEM_data[67]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__3_ ( .D(n2686), .CLK(clk), .Q(
        inst_data_MEM_data[35]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__3_ ( .D(n2654), .CLK(clk), .Q(
        inst_data_MEM_data[3]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__3_ ( .D(n2621), .CLK(clk), .Q(
        inst_data_MEM_data[195]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__3_ ( .D(n2615), .CLK(clk), .Q(
        inst_data_MEM_data[163]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__3_ ( .D(n2583), .CLK(clk), .Q(
        inst_data_MEM_data[131]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__3_ ( .D(n2554), .CLK(clk), .Q(
        inst_data_MEM_data[99]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__3_ ( .D(n2522), .CLK(clk), .Q(
        inst_data_MEM_data[227]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_3_ ( .D(inst_ID2EX_reg_N42), .CLK(clk), .Q(reg_read_data_1_EX[3]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_3_ ( .D(inst_EX2MEM_reg_N42), .CLK(
        clk), .Q(alu_result_MEM[3]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_3_ ( .D(u_MEM2WB_reg_N42), .CLK(clk), 
        .Q(alu_result_WB[3]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_4_ ( .D(u_MEM2WB_reg_N11), .CLK(clk), 
        .Q(mem_read_data_WB[4]) );
  DFFPOSX1 inst_register_registers_reg_7__4_ ( .D(n2465), .CLK(clk), .Q(
        inst_register_registers[228]) );
  DFFPOSX1 inst_register_registers_reg_6__4_ ( .D(n2408), .CLK(clk), .Q(
        inst_register_registers[196]) );
  DFFPOSX1 inst_register_registers_reg_5__4_ ( .D(n2402), .CLK(clk), .Q(
        inst_register_registers[164]) );
  DFFPOSX1 inst_register_registers_reg_4__4_ ( .D(n2370), .CLK(clk), .Q(
        inst_register_registers[132]) );
  DFFPOSX1 inst_register_registers_reg_3__4_ ( .D(n2341), .CLK(clk), .Q(
        inst_register_registers[100]) );
  DFFPOSX1 inst_register_registers_reg_2__4_ ( .D(n2305), .CLK(clk), .Q(
        inst_register_registers[68]) );
  DFFPOSX1 inst_register_registers_reg_1__4_ ( .D(n2273), .CLK(clk), .Q(
        inst_register_registers[36]) );
  DFFPOSX1 inst_register_registers_reg_0__4_ ( .D(n2241), .CLK(clk), .Q(
        inst_register_registers[4]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_4_ ( .D(inst_ID2EX_reg_N75), .CLK(clk), .Q(reg_read_data_2_EX[4]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_4_ ( .D(inst_EX2MEM_reg_N75), 
        .CLK(clk), .Q(write_mem_data_MEM[4]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__4_ ( .D(n2717), .CLK(clk), .Q(
        inst_data_MEM_data[68]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__4_ ( .D(n2685), .CLK(clk), .Q(
        inst_data_MEM_data[36]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__4_ ( .D(n2653), .CLK(clk), .Q(
        inst_data_MEM_data[4]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__4_ ( .D(n2620), .CLK(clk), .Q(
        inst_data_MEM_data[196]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__4_ ( .D(n2614), .CLK(clk), .Q(
        inst_data_MEM_data[164]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__4_ ( .D(n2582), .CLK(clk), .Q(
        inst_data_MEM_data[132]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__4_ ( .D(n2553), .CLK(clk), .Q(
        inst_data_MEM_data[100]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__4_ ( .D(n2521), .CLK(clk), .Q(
        inst_data_MEM_data[228]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_4_ ( .D(inst_ID2EX_reg_N43), .CLK(clk), .Q(reg_read_data_1_EX[4]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_4_ ( .D(inst_EX2MEM_reg_N43), .CLK(
        clk), .Q(alu_result_MEM[4]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_4_ ( .D(u_MEM2WB_reg_N43), .CLK(clk), 
        .Q(alu_result_WB[4]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_5_ ( .D(u_MEM2WB_reg_N12), .CLK(clk), 
        .Q(mem_read_data_WB[5]) );
  DFFPOSX1 inst_register_registers_reg_7__5_ ( .D(n2464), .CLK(clk), .Q(
        inst_register_registers[229]) );
  DFFPOSX1 inst_register_registers_reg_6__5_ ( .D(n2413), .CLK(clk), .Q(
        inst_register_registers[197]) );
  DFFPOSX1 inst_register_registers_reg_5__5_ ( .D(n2401), .CLK(clk), .Q(
        inst_register_registers[165]) );
  DFFPOSX1 inst_register_registers_reg_4__5_ ( .D(n2369), .CLK(clk), .Q(
        inst_register_registers[133]) );
  DFFPOSX1 inst_register_registers_reg_3__5_ ( .D(n2340), .CLK(clk), .Q(
        inst_register_registers[101]) );
  DFFPOSX1 inst_register_registers_reg_2__5_ ( .D(n2304), .CLK(clk), .Q(
        inst_register_registers[69]) );
  DFFPOSX1 inst_register_registers_reg_1__5_ ( .D(n2272), .CLK(clk), .Q(
        inst_register_registers[37]) );
  DFFPOSX1 inst_register_registers_reg_0__5_ ( .D(n2240), .CLK(clk), .Q(
        inst_register_registers[5]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_5_ ( .D(inst_ID2EX_reg_N76), .CLK(clk), .Q(reg_read_data_2_EX[5]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_5_ ( .D(inst_EX2MEM_reg_N76), 
        .CLK(clk), .Q(write_mem_data_MEM[5]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__5_ ( .D(n2716), .CLK(clk), .Q(
        inst_data_MEM_data[69]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__5_ ( .D(n2684), .CLK(clk), .Q(
        inst_data_MEM_data[37]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__5_ ( .D(n2652), .CLK(clk), .Q(
        inst_data_MEM_data[5]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__5_ ( .D(n2625), .CLK(clk), .Q(
        inst_data_MEM_data[197]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__5_ ( .D(n2613), .CLK(clk), .Q(
        inst_data_MEM_data[165]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__5_ ( .D(n2581), .CLK(clk), .Q(
        inst_data_MEM_data[133]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__5_ ( .D(n2552), .CLK(clk), .Q(
        inst_data_MEM_data[101]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__5_ ( .D(n2520), .CLK(clk), .Q(
        inst_data_MEM_data[229]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_5_ ( .D(inst_ID2EX_reg_N44), .CLK(clk), .Q(reg_read_data_1_EX[5]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_5_ ( .D(inst_EX2MEM_reg_N44), .CLK(
        clk), .Q(alu_result_MEM[5]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_5_ ( .D(u_MEM2WB_reg_N44), .CLK(clk), 
        .Q(alu_result_WB[5]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_6_ ( .D(u_MEM2WB_reg_N13), .CLK(clk), 
        .Q(mem_read_data_WB[6]) );
  DFFPOSX1 inst_register_registers_reg_7__6_ ( .D(n2463), .CLK(clk), .Q(
        inst_register_registers[230]) );
  DFFPOSX1 inst_register_registers_reg_6__6_ ( .D(n2439), .CLK(clk), .Q(
        inst_register_registers[198]) );
  DFFPOSX1 inst_register_registers_reg_5__6_ ( .D(n2400), .CLK(clk), .Q(
        inst_register_registers[166]) );
  DFFPOSX1 inst_register_registers_reg_4__6_ ( .D(n2368), .CLK(clk), .Q(
        inst_register_registers[134]) );
  DFFPOSX1 inst_register_registers_reg_3__6_ ( .D(n2339), .CLK(clk), .Q(
        inst_register_registers[102]) );
  DFFPOSX1 inst_register_registers_reg_2__6_ ( .D(n2303), .CLK(clk), .Q(
        inst_register_registers[70]) );
  DFFPOSX1 inst_register_registers_reg_1__6_ ( .D(n2271), .CLK(clk), .Q(
        inst_register_registers[38]) );
  DFFPOSX1 inst_register_registers_reg_0__6_ ( .D(n2239), .CLK(clk), .Q(
        inst_register_registers[6]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_6_ ( .D(inst_ID2EX_reg_N77), .CLK(clk), .Q(reg_read_data_2_EX[6]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_6_ ( .D(inst_EX2MEM_reg_N77), 
        .CLK(clk), .Q(write_mem_data_MEM[6]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__6_ ( .D(n2715), .CLK(clk), .Q(
        inst_data_MEM_data[70]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__6_ ( .D(n2683), .CLK(clk), .Q(
        inst_data_MEM_data[38]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__6_ ( .D(n2651), .CLK(clk), .Q(
        inst_data_MEM_data[6]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__6_ ( .D(n2612), .CLK(clk), .Q(
        inst_data_MEM_data[166]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__6_ ( .D(n2580), .CLK(clk), .Q(
        inst_data_MEM_data[134]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__6_ ( .D(n2551), .CLK(clk), .Q(
        inst_data_MEM_data[102]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__6_ ( .D(n2519), .CLK(clk), .Q(
        inst_data_MEM_data[230]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__6_ ( .D(n2495), .CLK(clk), .Q(
        inst_data_MEM_data[198]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_6_ ( .D(inst_ID2EX_reg_N45), .CLK(clk), .Q(reg_read_data_1_EX[6]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_6_ ( .D(inst_EX2MEM_reg_N45), .CLK(
        clk), .Q(alu_result_MEM[6]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_6_ ( .D(u_MEM2WB_reg_N45), .CLK(clk), 
        .Q(alu_result_WB[6]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_7_ ( .D(u_MEM2WB_reg_N14), .CLK(clk), 
        .Q(mem_read_data_WB[7]) );
  DFFPOSX1 inst_register_registers_reg_7__7_ ( .D(n2462), .CLK(clk), .Q(
        inst_register_registers[231]) );
  DFFPOSX1 inst_register_registers_reg_6__7_ ( .D(n2438), .CLK(clk), .Q(
        inst_register_registers[199]) );
  DFFPOSX1 inst_register_registers_reg_5__7_ ( .D(n2399), .CLK(clk), .Q(
        inst_register_registers[167]) );
  DFFPOSX1 inst_register_registers_reg_4__7_ ( .D(n2367), .CLK(clk), .Q(
        inst_register_registers[135]) );
  DFFPOSX1 inst_register_registers_reg_3__7_ ( .D(n2338), .CLK(clk), .Q(
        inst_register_registers[103]) );
  DFFPOSX1 inst_register_registers_reg_2__7_ ( .D(n2302), .CLK(clk), .Q(
        inst_register_registers[71]) );
  DFFPOSX1 inst_register_registers_reg_1__7_ ( .D(n2270), .CLK(clk), .Q(
        inst_register_registers[39]) );
  DFFPOSX1 inst_register_registers_reg_0__7_ ( .D(n2238), .CLK(clk), .Q(
        inst_register_registers[7]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_7_ ( .D(inst_ID2EX_reg_N78), .CLK(clk), .Q(reg_read_data_2_EX[7]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_7_ ( .D(inst_EX2MEM_reg_N78), 
        .CLK(clk), .Q(write_mem_data_MEM[7]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__7_ ( .D(n2714), .CLK(clk), .Q(
        inst_data_MEM_data[71]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__7_ ( .D(n2682), .CLK(clk), .Q(
        inst_data_MEM_data[39]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__7_ ( .D(n2650), .CLK(clk), .Q(
        inst_data_MEM_data[7]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__7_ ( .D(n2611), .CLK(clk), .Q(
        inst_data_MEM_data[167]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__7_ ( .D(n2579), .CLK(clk), .Q(
        inst_data_MEM_data[135]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__7_ ( .D(n2550), .CLK(clk), .Q(
        inst_data_MEM_data[103]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__7_ ( .D(n2518), .CLK(clk), .Q(
        inst_data_MEM_data[231]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__7_ ( .D(n2494), .CLK(clk), .Q(
        inst_data_MEM_data[199]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_7_ ( .D(inst_ID2EX_reg_N46), .CLK(clk), .Q(reg_read_data_1_EX[7]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_7_ ( .D(inst_EX2MEM_reg_N46), .CLK(
        clk), .Q(alu_result_MEM[7]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_7_ ( .D(u_MEM2WB_reg_N46), .CLK(clk), 
        .Q(alu_result_WB[7]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_8_ ( .D(u_MEM2WB_reg_N15), .CLK(clk), 
        .Q(mem_read_data_WB[8]) );
  DFFPOSX1 inst_register_registers_reg_7__8_ ( .D(n2461), .CLK(clk), .Q(
        inst_register_registers[232]) );
  DFFPOSX1 inst_register_registers_reg_6__8_ ( .D(n2437), .CLK(clk), .Q(
        inst_register_registers[200]) );
  DFFPOSX1 inst_register_registers_reg_5__8_ ( .D(n2398), .CLK(clk), .Q(
        inst_register_registers[168]) );
  DFFPOSX1 inst_register_registers_reg_4__8_ ( .D(n2366), .CLK(clk), .Q(
        inst_register_registers[136]) );
  DFFPOSX1 inst_register_registers_reg_3__8_ ( .D(n2337), .CLK(clk), .Q(
        inst_register_registers[104]) );
  DFFPOSX1 inst_register_registers_reg_2__8_ ( .D(n2301), .CLK(clk), .Q(
        inst_register_registers[72]) );
  DFFPOSX1 inst_register_registers_reg_1__8_ ( .D(n2269), .CLK(clk), .Q(
        inst_register_registers[40]) );
  DFFPOSX1 inst_register_registers_reg_0__8_ ( .D(n2237), .CLK(clk), .Q(
        inst_register_registers[8]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_8_ ( .D(inst_ID2EX_reg_N79), .CLK(clk), .Q(reg_read_data_2_EX[8]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_8_ ( .D(inst_EX2MEM_reg_N79), 
        .CLK(clk), .Q(write_mem_data_MEM[8]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__8_ ( .D(n2713), .CLK(clk), .Q(
        inst_data_MEM_data[72]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__8_ ( .D(n2681), .CLK(clk), .Q(
        inst_data_MEM_data[40]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__8_ ( .D(n2649), .CLK(clk), .Q(
        inst_data_MEM_data[8]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__8_ ( .D(n2610), .CLK(clk), .Q(
        inst_data_MEM_data[168]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__8_ ( .D(n2578), .CLK(clk), .Q(
        inst_data_MEM_data[136]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__8_ ( .D(n2549), .CLK(clk), .Q(
        inst_data_MEM_data[104]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__8_ ( .D(n2517), .CLK(clk), .Q(
        inst_data_MEM_data[232]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__8_ ( .D(n2493), .CLK(clk), .Q(
        inst_data_MEM_data[200]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_8_ ( .D(inst_ID2EX_reg_N47), .CLK(clk), .Q(reg_read_data_1_EX[8]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_8_ ( .D(inst_EX2MEM_reg_N47), .CLK(
        clk), .Q(alu_result_MEM[8]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_8_ ( .D(u_MEM2WB_reg_N47), .CLK(clk), 
        .Q(alu_result_WB[8]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_9_ ( .D(u_MEM2WB_reg_N16), .CLK(clk), 
        .Q(mem_read_data_WB[9]) );
  DFFPOSX1 inst_register_registers_reg_7__9_ ( .D(n2460), .CLK(clk), .Q(
        inst_register_registers[233]) );
  DFFPOSX1 inst_register_registers_reg_6__9_ ( .D(n2436), .CLK(clk), .Q(
        inst_register_registers[201]) );
  DFFPOSX1 inst_register_registers_reg_5__9_ ( .D(n2397), .CLK(clk), .Q(
        inst_register_registers[169]) );
  DFFPOSX1 inst_register_registers_reg_4__9_ ( .D(n2365), .CLK(clk), .Q(
        inst_register_registers[137]) );
  DFFPOSX1 inst_register_registers_reg_3__9_ ( .D(n2336), .CLK(clk), .Q(
        inst_register_registers[105]) );
  DFFPOSX1 inst_register_registers_reg_2__9_ ( .D(n2300), .CLK(clk), .Q(
        inst_register_registers[73]) );
  DFFPOSX1 inst_register_registers_reg_1__9_ ( .D(n2268), .CLK(clk), .Q(
        inst_register_registers[41]) );
  DFFPOSX1 inst_register_registers_reg_0__9_ ( .D(n2236), .CLK(clk), .Q(
        inst_register_registers[9]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_9_ ( .D(inst_ID2EX_reg_N80), .CLK(clk), .Q(reg_read_data_2_EX[9]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_9_ ( .D(inst_EX2MEM_reg_N80), 
        .CLK(clk), .Q(write_mem_data_MEM[9]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__9_ ( .D(n2712), .CLK(clk), .Q(
        inst_data_MEM_data[73]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__9_ ( .D(n2680), .CLK(clk), .Q(
        inst_data_MEM_data[41]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__9_ ( .D(n2648), .CLK(clk), .Q(
        inst_data_MEM_data[9]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__9_ ( .D(n2609), .CLK(clk), .Q(
        inst_data_MEM_data[169]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__9_ ( .D(n2577), .CLK(clk), .Q(
        inst_data_MEM_data[137]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__9_ ( .D(n2548), .CLK(clk), .Q(
        inst_data_MEM_data[105]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__9_ ( .D(n2516), .CLK(clk), .Q(
        inst_data_MEM_data[233]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__9_ ( .D(n2492), .CLK(clk), .Q(
        inst_data_MEM_data[201]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_9_ ( .D(inst_ID2EX_reg_N48), .CLK(clk), .Q(reg_read_data_1_EX[9]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_9_ ( .D(inst_EX2MEM_reg_N48), .CLK(
        clk), .Q(alu_result_MEM[9]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_9_ ( .D(u_MEM2WB_reg_N48), .CLK(clk), 
        .Q(alu_result_WB[9]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_10_ ( .D(u_MEM2WB_reg_N17), .CLK(clk), 
        .Q(mem_read_data_WB[10]) );
  DFFPOSX1 inst_register_registers_reg_7__10_ ( .D(n2459), .CLK(clk), .Q(
        inst_register_registers[234]) );
  DFFPOSX1 inst_register_registers_reg_6__10_ ( .D(n2435), .CLK(clk), .Q(
        inst_register_registers[202]) );
  DFFPOSX1 inst_register_registers_reg_5__10_ ( .D(n2396), .CLK(clk), .Q(
        inst_register_registers[170]) );
  DFFPOSX1 inst_register_registers_reg_4__10_ ( .D(n2364), .CLK(clk), .Q(
        inst_register_registers[138]) );
  DFFPOSX1 inst_register_registers_reg_3__10_ ( .D(n2335), .CLK(clk), .Q(
        inst_register_registers[106]) );
  DFFPOSX1 inst_register_registers_reg_2__10_ ( .D(n2299), .CLK(clk), .Q(
        inst_register_registers[74]) );
  DFFPOSX1 inst_register_registers_reg_1__10_ ( .D(n2267), .CLK(clk), .Q(
        inst_register_registers[42]) );
  DFFPOSX1 inst_register_registers_reg_0__10_ ( .D(n2235), .CLK(clk), .Q(
        inst_register_registers[10]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_10_ ( .D(inst_ID2EX_reg_N81), .CLK(
        clk), .Q(reg_read_data_2_EX[10]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_10_ ( .D(inst_EX2MEM_reg_N81), 
        .CLK(clk), .Q(write_mem_data_MEM[10]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__10_ ( .D(n2711), .CLK(clk), .Q(
        inst_data_MEM_data[74]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__10_ ( .D(n2679), .CLK(clk), .Q(
        inst_data_MEM_data[42]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__10_ ( .D(n2647), .CLK(clk), .Q(
        inst_data_MEM_data[10]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__10_ ( .D(n2608), .CLK(clk), .Q(
        inst_data_MEM_data[170]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__10_ ( .D(n2576), .CLK(clk), .Q(
        inst_data_MEM_data[138]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__10_ ( .D(n2547), .CLK(clk), .Q(
        inst_data_MEM_data[106]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__10_ ( .D(n2515), .CLK(clk), .Q(
        inst_data_MEM_data[234]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__10_ ( .D(n2491), .CLK(clk), .Q(
        inst_data_MEM_data[202]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_10_ ( .D(inst_ID2EX_reg_N49), .CLK(
        clk), .Q(reg_read_data_1_EX[10]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_10_ ( .D(inst_EX2MEM_reg_N49), .CLK(
        clk), .Q(alu_result_MEM[10]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_10_ ( .D(u_MEM2WB_reg_N49), .CLK(clk), 
        .Q(alu_result_WB[10]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_11_ ( .D(u_MEM2WB_reg_N18), .CLK(clk), 
        .Q(mem_read_data_WB[11]) );
  DFFPOSX1 inst_register_registers_reg_7__11_ ( .D(n2458), .CLK(clk), .Q(
        inst_register_registers[235]) );
  DFFPOSX1 inst_register_registers_reg_6__11_ ( .D(n2434), .CLK(clk), .Q(
        inst_register_registers[203]) );
  DFFPOSX1 inst_register_registers_reg_5__11_ ( .D(n2395), .CLK(clk), .Q(
        inst_register_registers[171]) );
  DFFPOSX1 inst_register_registers_reg_4__11_ ( .D(n2363), .CLK(clk), .Q(
        inst_register_registers[139]) );
  DFFPOSX1 inst_register_registers_reg_3__11_ ( .D(n2334), .CLK(clk), .Q(
        inst_register_registers[107]) );
  DFFPOSX1 inst_register_registers_reg_2__11_ ( .D(n2298), .CLK(clk), .Q(
        inst_register_registers[75]) );
  DFFPOSX1 inst_register_registers_reg_1__11_ ( .D(n2266), .CLK(clk), .Q(
        inst_register_registers[43]) );
  DFFPOSX1 inst_register_registers_reg_0__11_ ( .D(n2234), .CLK(clk), .Q(
        inst_register_registers[11]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_11_ ( .D(inst_ID2EX_reg_N82), .CLK(
        clk), .Q(reg_read_data_2_EX[11]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_11_ ( .D(inst_EX2MEM_reg_N82), 
        .CLK(clk), .Q(write_mem_data_MEM[11]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__11_ ( .D(n2710), .CLK(clk), .Q(
        inst_data_MEM_data[75]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__11_ ( .D(n2678), .CLK(clk), .Q(
        inst_data_MEM_data[43]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__11_ ( .D(n2646), .CLK(clk), .Q(
        inst_data_MEM_data[11]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__11_ ( .D(n2607), .CLK(clk), .Q(
        inst_data_MEM_data[171]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__11_ ( .D(n2575), .CLK(clk), .Q(
        inst_data_MEM_data[139]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__11_ ( .D(n2546), .CLK(clk), .Q(
        inst_data_MEM_data[107]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__11_ ( .D(n2514), .CLK(clk), .Q(
        inst_data_MEM_data[235]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__11_ ( .D(n2490), .CLK(clk), .Q(
        inst_data_MEM_data[203]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_11_ ( .D(inst_ID2EX_reg_N50), .CLK(
        clk), .Q(reg_read_data_1_EX[11]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_11_ ( .D(inst_EX2MEM_reg_N50), .CLK(
        clk), .Q(alu_result_MEM[11]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_11_ ( .D(u_MEM2WB_reg_N50), .CLK(clk), 
        .Q(alu_result_WB[11]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_12_ ( .D(u_MEM2WB_reg_N19), .CLK(clk), 
        .Q(mem_read_data_WB[12]) );
  DFFPOSX1 inst_register_registers_reg_7__12_ ( .D(n2457), .CLK(clk), .Q(
        inst_register_registers[236]) );
  DFFPOSX1 inst_register_registers_reg_6__12_ ( .D(n2433), .CLK(clk), .Q(
        inst_register_registers[204]) );
  DFFPOSX1 inst_register_registers_reg_5__12_ ( .D(n2394), .CLK(clk), .Q(
        inst_register_registers[172]) );
  DFFPOSX1 inst_register_registers_reg_4__12_ ( .D(n2362), .CLK(clk), .Q(
        inst_register_registers[140]) );
  DFFPOSX1 inst_register_registers_reg_3__12_ ( .D(n2333), .CLK(clk), .Q(
        inst_register_registers[108]) );
  DFFPOSX1 inst_register_registers_reg_2__12_ ( .D(n2297), .CLK(clk), .Q(
        inst_register_registers[76]) );
  DFFPOSX1 inst_register_registers_reg_1__12_ ( .D(n2265), .CLK(clk), .Q(
        inst_register_registers[44]) );
  DFFPOSX1 inst_register_registers_reg_0__12_ ( .D(n2233), .CLK(clk), .Q(
        inst_register_registers[12]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_12_ ( .D(inst_ID2EX_reg_N83), .CLK(
        clk), .Q(reg_read_data_2_EX[12]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_12_ ( .D(inst_EX2MEM_reg_N83), 
        .CLK(clk), .Q(write_mem_data_MEM[12]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__12_ ( .D(n2709), .CLK(clk), .Q(
        inst_data_MEM_data[76]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__12_ ( .D(n2677), .CLK(clk), .Q(
        inst_data_MEM_data[44]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__12_ ( .D(n2645), .CLK(clk), .Q(
        inst_data_MEM_data[12]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__12_ ( .D(n2606), .CLK(clk), .Q(
        inst_data_MEM_data[172]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__12_ ( .D(n2574), .CLK(clk), .Q(
        inst_data_MEM_data[140]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__12_ ( .D(n2545), .CLK(clk), .Q(
        inst_data_MEM_data[108]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__12_ ( .D(n2513), .CLK(clk), .Q(
        inst_data_MEM_data[236]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__12_ ( .D(n2489), .CLK(clk), .Q(
        inst_data_MEM_data[204]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_12_ ( .D(inst_ID2EX_reg_N51), .CLK(
        clk), .Q(reg_read_data_1_EX[12]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_12_ ( .D(inst_EX2MEM_reg_N51), .CLK(
        clk), .Q(alu_result_MEM[12]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_12_ ( .D(u_MEM2WB_reg_N51), .CLK(clk), 
        .Q(alu_result_WB[12]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_13_ ( .D(u_MEM2WB_reg_N20), .CLK(clk), 
        .Q(mem_read_data_WB[13]) );
  DFFPOSX1 inst_register_registers_reg_7__13_ ( .D(n2456), .CLK(clk), .Q(
        inst_register_registers[237]) );
  DFFPOSX1 inst_register_registers_reg_6__13_ ( .D(n2432), .CLK(clk), .Q(
        inst_register_registers[205]) );
  DFFPOSX1 inst_register_registers_reg_5__13_ ( .D(n2393), .CLK(clk), .Q(
        inst_register_registers[173]) );
  DFFPOSX1 inst_register_registers_reg_4__13_ ( .D(n2361), .CLK(clk), .Q(
        inst_register_registers[141]) );
  DFFPOSX1 inst_register_registers_reg_3__13_ ( .D(n2332), .CLK(clk), .Q(
        inst_register_registers[109]) );
  DFFPOSX1 inst_register_registers_reg_2__13_ ( .D(n2296), .CLK(clk), .Q(
        inst_register_registers[77]) );
  DFFPOSX1 inst_register_registers_reg_1__13_ ( .D(n2264), .CLK(clk), .Q(
        inst_register_registers[45]) );
  DFFPOSX1 inst_register_registers_reg_0__13_ ( .D(n2232), .CLK(clk), .Q(
        inst_register_registers[13]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_13_ ( .D(inst_ID2EX_reg_N84), .CLK(
        clk), .Q(reg_read_data_2_EX[13]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_13_ ( .D(inst_EX2MEM_reg_N84), 
        .CLK(clk), .Q(write_mem_data_MEM[13]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__13_ ( .D(n2708), .CLK(clk), .Q(
        inst_data_MEM_data[77]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__13_ ( .D(n2676), .CLK(clk), .Q(
        inst_data_MEM_data[45]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__13_ ( .D(n2644), .CLK(clk), .Q(
        inst_data_MEM_data[13]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__13_ ( .D(n2605), .CLK(clk), .Q(
        inst_data_MEM_data[173]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__13_ ( .D(n2573), .CLK(clk), .Q(
        inst_data_MEM_data[141]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__13_ ( .D(n2544), .CLK(clk), .Q(
        inst_data_MEM_data[109]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__13_ ( .D(n2512), .CLK(clk), .Q(
        inst_data_MEM_data[237]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__13_ ( .D(n2488), .CLK(clk), .Q(
        inst_data_MEM_data[205]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_13_ ( .D(inst_ID2EX_reg_N52), .CLK(
        clk), .Q(reg_read_data_1_EX[13]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_13_ ( .D(inst_EX2MEM_reg_N52), .CLK(
        clk), .Q(alu_result_MEM[13]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_13_ ( .D(u_MEM2WB_reg_N52), .CLK(clk), 
        .Q(alu_result_WB[13]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_14_ ( .D(u_MEM2WB_reg_N21), .CLK(clk), 
        .Q(mem_read_data_WB[14]) );
  DFFPOSX1 inst_register_registers_reg_7__14_ ( .D(n2455), .CLK(clk), .Q(
        inst_register_registers[238]) );
  DFFPOSX1 inst_register_registers_reg_6__14_ ( .D(n2431), .CLK(clk), .Q(
        inst_register_registers[206]) );
  DFFPOSX1 inst_register_registers_reg_5__14_ ( .D(n2392), .CLK(clk), .Q(
        inst_register_registers[174]) );
  DFFPOSX1 inst_register_registers_reg_4__14_ ( .D(n2360), .CLK(clk), .Q(
        inst_register_registers[142]) );
  DFFPOSX1 inst_register_registers_reg_3__14_ ( .D(n2331), .CLK(clk), .Q(
        inst_register_registers[110]) );
  DFFPOSX1 inst_register_registers_reg_2__14_ ( .D(n2295), .CLK(clk), .Q(
        inst_register_registers[78]) );
  DFFPOSX1 inst_register_registers_reg_1__14_ ( .D(n2263), .CLK(clk), .Q(
        inst_register_registers[46]) );
  DFFPOSX1 inst_register_registers_reg_0__14_ ( .D(n2231), .CLK(clk), .Q(
        inst_register_registers[14]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_14_ ( .D(inst_ID2EX_reg_N85), .CLK(
        clk), .Q(reg_read_data_2_EX[14]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_14_ ( .D(inst_EX2MEM_reg_N85), 
        .CLK(clk), .Q(write_mem_data_MEM[14]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__14_ ( .D(n2707), .CLK(clk), .Q(
        inst_data_MEM_data[78]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__14_ ( .D(n2675), .CLK(clk), .Q(
        inst_data_MEM_data[46]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__14_ ( .D(n2643), .CLK(clk), .Q(
        inst_data_MEM_data[14]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__14_ ( .D(n2604), .CLK(clk), .Q(
        inst_data_MEM_data[174]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__14_ ( .D(n2572), .CLK(clk), .Q(
        inst_data_MEM_data[142]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__14_ ( .D(n2543), .CLK(clk), .Q(
        inst_data_MEM_data[110]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__14_ ( .D(n2511), .CLK(clk), .Q(
        inst_data_MEM_data[238]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__14_ ( .D(n2487), .CLK(clk), .Q(
        inst_data_MEM_data[206]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_14_ ( .D(inst_ID2EX_reg_N53), .CLK(
        clk), .Q(reg_read_data_1_EX[14]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_14_ ( .D(inst_EX2MEM_reg_N53), .CLK(
        clk), .Q(alu_result_MEM[14]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_14_ ( .D(u_MEM2WB_reg_N53), .CLK(clk), 
        .Q(alu_result_WB[14]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_15_ ( .D(u_MEM2WB_reg_N22), .CLK(clk), 
        .Q(mem_read_data_WB[15]) );
  DFFPOSX1 inst_register_registers_reg_7__15_ ( .D(n2454), .CLK(clk), .Q(
        inst_register_registers[239]) );
  DFFPOSX1 inst_register_registers_reg_6__15_ ( .D(n2430), .CLK(clk), .Q(
        inst_register_registers[207]) );
  DFFPOSX1 inst_register_registers_reg_5__15_ ( .D(n2391), .CLK(clk), .Q(
        inst_register_registers[175]) );
  DFFPOSX1 inst_register_registers_reg_4__15_ ( .D(n2359), .CLK(clk), .Q(
        inst_register_registers[143]) );
  DFFPOSX1 inst_register_registers_reg_3__15_ ( .D(n2330), .CLK(clk), .Q(
        inst_register_registers[111]) );
  DFFPOSX1 inst_register_registers_reg_2__15_ ( .D(n2294), .CLK(clk), .Q(
        inst_register_registers[79]) );
  DFFPOSX1 inst_register_registers_reg_1__15_ ( .D(n2262), .CLK(clk), .Q(
        inst_register_registers[47]) );
  DFFPOSX1 inst_register_registers_reg_0__15_ ( .D(n2230), .CLK(clk), .Q(
        inst_register_registers[15]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_15_ ( .D(inst_ID2EX_reg_N86), .CLK(
        clk), .Q(reg_read_data_2_EX[15]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_15_ ( .D(inst_EX2MEM_reg_N86), 
        .CLK(clk), .Q(write_mem_data_MEM[15]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__15_ ( .D(n2706), .CLK(clk), .Q(
        inst_data_MEM_data[79]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__15_ ( .D(n2674), .CLK(clk), .Q(
        inst_data_MEM_data[47]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__15_ ( .D(n2642), .CLK(clk), .Q(
        inst_data_MEM_data[15]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__15_ ( .D(n2603), .CLK(clk), .Q(
        inst_data_MEM_data[175]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__15_ ( .D(n2571), .CLK(clk), .Q(
        inst_data_MEM_data[143]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__15_ ( .D(n2542), .CLK(clk), .Q(
        inst_data_MEM_data[111]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__15_ ( .D(n2510), .CLK(clk), .Q(
        inst_data_MEM_data[239]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__15_ ( .D(n2486), .CLK(clk), .Q(
        inst_data_MEM_data[207]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_15_ ( .D(inst_ID2EX_reg_N54), .CLK(
        clk), .Q(reg_read_data_1_EX[15]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_15_ ( .D(inst_EX2MEM_reg_N54), .CLK(
        clk), .Q(alu_result_MEM[15]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_15_ ( .D(u_MEM2WB_reg_N54), .CLK(clk), 
        .Q(alu_result_WB[15]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_16_ ( .D(u_MEM2WB_reg_N23), .CLK(clk), 
        .Q(mem_read_data_WB[16]) );
  DFFPOSX1 inst_register_registers_reg_7__16_ ( .D(n2453), .CLK(clk), .Q(
        inst_register_registers[240]) );
  DFFPOSX1 inst_register_registers_reg_6__16_ ( .D(n2429), .CLK(clk), .Q(
        inst_register_registers[208]) );
  DFFPOSX1 inst_register_registers_reg_5__16_ ( .D(n2390), .CLK(clk), .Q(
        inst_register_registers[176]) );
  DFFPOSX1 inst_register_registers_reg_4__16_ ( .D(n2358), .CLK(clk), .Q(
        inst_register_registers[144]) );
  DFFPOSX1 inst_register_registers_reg_3__16_ ( .D(n2329), .CLK(clk), .Q(
        inst_register_registers[112]) );
  DFFPOSX1 inst_register_registers_reg_2__16_ ( .D(n2293), .CLK(clk), .Q(
        inst_register_registers[80]) );
  DFFPOSX1 inst_register_registers_reg_1__16_ ( .D(n2261), .CLK(clk), .Q(
        inst_register_registers[48]) );
  DFFPOSX1 inst_register_registers_reg_0__16_ ( .D(n2229), .CLK(clk), .Q(
        inst_register_registers[16]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_16_ ( .D(inst_ID2EX_reg_N87), .CLK(
        clk), .Q(reg_read_data_2_EX[16]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_16_ ( .D(inst_EX2MEM_reg_N87), 
        .CLK(clk), .Q(write_mem_data_MEM[16]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__16_ ( .D(n2705), .CLK(clk), .Q(
        inst_data_MEM_data[80]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__16_ ( .D(n2673), .CLK(clk), .Q(
        inst_data_MEM_data[48]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__16_ ( .D(n2641), .CLK(clk), .Q(
        inst_data_MEM_data[16]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__16_ ( .D(n2602), .CLK(clk), .Q(
        inst_data_MEM_data[176]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__16_ ( .D(n2570), .CLK(clk), .Q(
        inst_data_MEM_data[144]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__16_ ( .D(n2541), .CLK(clk), .Q(
        inst_data_MEM_data[112]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__16_ ( .D(n2509), .CLK(clk), .Q(
        inst_data_MEM_data[240]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__16_ ( .D(n2485), .CLK(clk), .Q(
        inst_data_MEM_data[208]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_16_ ( .D(inst_ID2EX_reg_N55), .CLK(
        clk), .Q(reg_read_data_1_EX[16]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_16_ ( .D(inst_EX2MEM_reg_N55), .CLK(
        clk), .Q(alu_result_MEM[16]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_16_ ( .D(u_MEM2WB_reg_N55), .CLK(clk), 
        .Q(alu_result_WB[16]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_17_ ( .D(u_MEM2WB_reg_N24), .CLK(clk), 
        .Q(mem_read_data_WB[17]) );
  DFFPOSX1 inst_register_registers_reg_7__17_ ( .D(n2452), .CLK(clk), .Q(
        inst_register_registers[241]) );
  DFFPOSX1 inst_register_registers_reg_6__17_ ( .D(n2428), .CLK(clk), .Q(
        inst_register_registers[209]) );
  DFFPOSX1 inst_register_registers_reg_5__17_ ( .D(n2389), .CLK(clk), .Q(
        inst_register_registers[177]) );
  DFFPOSX1 inst_register_registers_reg_4__17_ ( .D(n2357), .CLK(clk), .Q(
        inst_register_registers[145]) );
  DFFPOSX1 inst_register_registers_reg_3__17_ ( .D(n2328), .CLK(clk), .Q(
        inst_register_registers[113]) );
  DFFPOSX1 inst_register_registers_reg_2__17_ ( .D(n2292), .CLK(clk), .Q(
        inst_register_registers[81]) );
  DFFPOSX1 inst_register_registers_reg_1__17_ ( .D(n2260), .CLK(clk), .Q(
        inst_register_registers[49]) );
  DFFPOSX1 inst_register_registers_reg_0__17_ ( .D(n2228), .CLK(clk), .Q(
        inst_register_registers[17]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_17_ ( .D(inst_ID2EX_reg_N88), .CLK(
        clk), .Q(reg_read_data_2_EX[17]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_17_ ( .D(inst_EX2MEM_reg_N88), 
        .CLK(clk), .Q(write_mem_data_MEM[17]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__17_ ( .D(n2704), .CLK(clk), .Q(
        inst_data_MEM_data[81]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__17_ ( .D(n2672), .CLK(clk), .Q(
        inst_data_MEM_data[49]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__17_ ( .D(n2640), .CLK(clk), .Q(
        inst_data_MEM_data[17]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__17_ ( .D(n2601), .CLK(clk), .Q(
        inst_data_MEM_data[177]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__17_ ( .D(n2569), .CLK(clk), .Q(
        inst_data_MEM_data[145]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__17_ ( .D(n2540), .CLK(clk), .Q(
        inst_data_MEM_data[113]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__17_ ( .D(n2508), .CLK(clk), .Q(
        inst_data_MEM_data[241]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__17_ ( .D(n2484), .CLK(clk), .Q(
        inst_data_MEM_data[209]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_17_ ( .D(inst_ID2EX_reg_N56), .CLK(
        clk), .Q(reg_read_data_1_EX[17]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_17_ ( .D(inst_EX2MEM_reg_N56), .CLK(
        clk), .Q(alu_result_MEM[17]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_17_ ( .D(u_MEM2WB_reg_N56), .CLK(clk), 
        .Q(alu_result_WB[17]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_18_ ( .D(u_MEM2WB_reg_N25), .CLK(clk), 
        .Q(mem_read_data_WB[18]) );
  DFFPOSX1 inst_register_registers_reg_7__18_ ( .D(n2451), .CLK(clk), .Q(
        inst_register_registers[242]) );
  DFFPOSX1 inst_register_registers_reg_6__18_ ( .D(n2427), .CLK(clk), .Q(
        inst_register_registers[210]) );
  DFFPOSX1 inst_register_registers_reg_5__18_ ( .D(n2388), .CLK(clk), .Q(
        inst_register_registers[178]) );
  DFFPOSX1 inst_register_registers_reg_4__18_ ( .D(n2356), .CLK(clk), .Q(
        inst_register_registers[146]) );
  DFFPOSX1 inst_register_registers_reg_3__18_ ( .D(n2327), .CLK(clk), .Q(
        inst_register_registers[114]) );
  DFFPOSX1 inst_register_registers_reg_2__18_ ( .D(n2291), .CLK(clk), .Q(
        inst_register_registers[82]) );
  DFFPOSX1 inst_register_registers_reg_1__18_ ( .D(n2259), .CLK(clk), .Q(
        inst_register_registers[50]) );
  DFFPOSX1 inst_register_registers_reg_0__18_ ( .D(n2227), .CLK(clk), .Q(
        inst_register_registers[18]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_18_ ( .D(inst_ID2EX_reg_N89), .CLK(
        clk), .Q(reg_read_data_2_EX[18]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_18_ ( .D(inst_EX2MEM_reg_N89), 
        .CLK(clk), .Q(write_mem_data_MEM[18]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__18_ ( .D(n2703), .CLK(clk), .Q(
        inst_data_MEM_data[82]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__18_ ( .D(n2671), .CLK(clk), .Q(
        inst_data_MEM_data[50]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__18_ ( .D(n2639), .CLK(clk), .Q(
        inst_data_MEM_data[18]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__18_ ( .D(n2600), .CLK(clk), .Q(
        inst_data_MEM_data[178]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__18_ ( .D(n2568), .CLK(clk), .Q(
        inst_data_MEM_data[146]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__18_ ( .D(n2539), .CLK(clk), .Q(
        inst_data_MEM_data[114]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__18_ ( .D(n2507), .CLK(clk), .Q(
        inst_data_MEM_data[242]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__18_ ( .D(n2483), .CLK(clk), .Q(
        inst_data_MEM_data[210]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_18_ ( .D(inst_ID2EX_reg_N57), .CLK(
        clk), .Q(reg_read_data_1_EX[18]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_18_ ( .D(inst_EX2MEM_reg_N57), .CLK(
        clk), .Q(alu_result_MEM[18]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_18_ ( .D(u_MEM2WB_reg_N57), .CLK(clk), 
        .Q(alu_result_WB[18]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_19_ ( .D(u_MEM2WB_reg_N26), .CLK(clk), 
        .Q(mem_read_data_WB[19]) );
  DFFPOSX1 inst_register_registers_reg_7__19_ ( .D(n2450), .CLK(clk), .Q(
        inst_register_registers[243]) );
  DFFPOSX1 inst_register_registers_reg_6__19_ ( .D(n2426), .CLK(clk), .Q(
        inst_register_registers[211]) );
  DFFPOSX1 inst_register_registers_reg_5__19_ ( .D(n2387), .CLK(clk), .Q(
        inst_register_registers[179]) );
  DFFPOSX1 inst_register_registers_reg_4__19_ ( .D(n2355), .CLK(clk), .Q(
        inst_register_registers[147]) );
  DFFPOSX1 inst_register_registers_reg_3__19_ ( .D(n2326), .CLK(clk), .Q(
        inst_register_registers[115]) );
  DFFPOSX1 inst_register_registers_reg_2__19_ ( .D(n2290), .CLK(clk), .Q(
        inst_register_registers[83]) );
  DFFPOSX1 inst_register_registers_reg_1__19_ ( .D(n2258), .CLK(clk), .Q(
        inst_register_registers[51]) );
  DFFPOSX1 inst_register_registers_reg_0__19_ ( .D(n2226), .CLK(clk), .Q(
        inst_register_registers[19]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_19_ ( .D(inst_ID2EX_reg_N90), .CLK(
        clk), .Q(reg_read_data_2_EX[19]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_19_ ( .D(inst_EX2MEM_reg_N90), 
        .CLK(clk), .Q(write_mem_data_MEM[19]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__19_ ( .D(n2702), .CLK(clk), .Q(
        inst_data_MEM_data[83]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__19_ ( .D(n2670), .CLK(clk), .Q(
        inst_data_MEM_data[51]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__19_ ( .D(n2638), .CLK(clk), .Q(
        inst_data_MEM_data[19]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__19_ ( .D(n2599), .CLK(clk), .Q(
        inst_data_MEM_data[179]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__19_ ( .D(n2567), .CLK(clk), .Q(
        inst_data_MEM_data[147]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__19_ ( .D(n2538), .CLK(clk), .Q(
        inst_data_MEM_data[115]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__19_ ( .D(n2506), .CLK(clk), .Q(
        inst_data_MEM_data[243]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__19_ ( .D(n2482), .CLK(clk), .Q(
        inst_data_MEM_data[211]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_19_ ( .D(inst_ID2EX_reg_N58), .CLK(
        clk), .Q(reg_read_data_1_EX[19]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_19_ ( .D(inst_EX2MEM_reg_N58), .CLK(
        clk), .Q(alu_result_MEM[19]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_19_ ( .D(u_MEM2WB_reg_N58), .CLK(clk), 
        .Q(alu_result_WB[19]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_20_ ( .D(u_MEM2WB_reg_N27), .CLK(clk), 
        .Q(mem_read_data_WB[20]) );
  DFFPOSX1 inst_register_registers_reg_7__20_ ( .D(n2449), .CLK(clk), .Q(
        inst_register_registers[244]) );
  DFFPOSX1 inst_register_registers_reg_6__20_ ( .D(n2425), .CLK(clk), .Q(
        inst_register_registers[212]) );
  DFFPOSX1 inst_register_registers_reg_5__20_ ( .D(n2386), .CLK(clk), .Q(
        inst_register_registers[180]) );
  DFFPOSX1 inst_register_registers_reg_4__20_ ( .D(n2354), .CLK(clk), .Q(
        inst_register_registers[148]) );
  DFFPOSX1 inst_register_registers_reg_3__20_ ( .D(n2325), .CLK(clk), .Q(
        inst_register_registers[116]) );
  DFFPOSX1 inst_register_registers_reg_2__20_ ( .D(n2289), .CLK(clk), .Q(
        inst_register_registers[84]) );
  DFFPOSX1 inst_register_registers_reg_1__20_ ( .D(n2257), .CLK(clk), .Q(
        inst_register_registers[52]) );
  DFFPOSX1 inst_register_registers_reg_0__20_ ( .D(n2225), .CLK(clk), .Q(
        inst_register_registers[20]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_20_ ( .D(inst_ID2EX_reg_N91), .CLK(
        clk), .Q(reg_read_data_2_EX[20]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_20_ ( .D(inst_EX2MEM_reg_N91), 
        .CLK(clk), .Q(write_mem_data_MEM[20]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__20_ ( .D(n2701), .CLK(clk), .Q(
        inst_data_MEM_data[84]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__20_ ( .D(n2669), .CLK(clk), .Q(
        inst_data_MEM_data[52]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__20_ ( .D(n2637), .CLK(clk), .Q(
        inst_data_MEM_data[20]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__20_ ( .D(n2598), .CLK(clk), .Q(
        inst_data_MEM_data[180]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__20_ ( .D(n2566), .CLK(clk), .Q(
        inst_data_MEM_data[148]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__20_ ( .D(n2537), .CLK(clk), .Q(
        inst_data_MEM_data[116]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__20_ ( .D(n2505), .CLK(clk), .Q(
        inst_data_MEM_data[244]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__20_ ( .D(n2481), .CLK(clk), .Q(
        inst_data_MEM_data[212]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_20_ ( .D(inst_ID2EX_reg_N59), .CLK(
        clk), .Q(reg_read_data_1_EX[20]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_20_ ( .D(inst_EX2MEM_reg_N59), .CLK(
        clk), .Q(alu_result_MEM[20]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_20_ ( .D(u_MEM2WB_reg_N59), .CLK(clk), 
        .Q(alu_result_WB[20]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_21_ ( .D(u_MEM2WB_reg_N28), .CLK(clk), 
        .Q(mem_read_data_WB[21]) );
  DFFPOSX1 inst_register_registers_reg_7__21_ ( .D(n2448), .CLK(clk), .Q(
        inst_register_registers[245]) );
  DFFPOSX1 inst_register_registers_reg_6__21_ ( .D(n2424), .CLK(clk), .Q(
        inst_register_registers[213]) );
  DFFPOSX1 inst_register_registers_reg_5__21_ ( .D(n2385), .CLK(clk), .Q(
        inst_register_registers[181]) );
  DFFPOSX1 inst_register_registers_reg_4__21_ ( .D(n2353), .CLK(clk), .Q(
        inst_register_registers[149]) );
  DFFPOSX1 inst_register_registers_reg_3__21_ ( .D(n2324), .CLK(clk), .Q(
        inst_register_registers[117]) );
  DFFPOSX1 inst_register_registers_reg_2__21_ ( .D(n2288), .CLK(clk), .Q(
        inst_register_registers[85]) );
  DFFPOSX1 inst_register_registers_reg_1__21_ ( .D(n2256), .CLK(clk), .Q(
        inst_register_registers[53]) );
  DFFPOSX1 inst_register_registers_reg_0__21_ ( .D(n2224), .CLK(clk), .Q(
        inst_register_registers[21]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_21_ ( .D(inst_ID2EX_reg_N92), .CLK(
        clk), .Q(reg_read_data_2_EX[21]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_21_ ( .D(inst_EX2MEM_reg_N92), 
        .CLK(clk), .Q(write_mem_data_MEM[21]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__21_ ( .D(n2700), .CLK(clk), .Q(
        inst_data_MEM_data[85]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__21_ ( .D(n2668), .CLK(clk), .Q(
        inst_data_MEM_data[53]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__21_ ( .D(n2636), .CLK(clk), .Q(
        inst_data_MEM_data[21]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__21_ ( .D(n2597), .CLK(clk), .Q(
        inst_data_MEM_data[181]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__21_ ( .D(n2565), .CLK(clk), .Q(
        inst_data_MEM_data[149]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__21_ ( .D(n2536), .CLK(clk), .Q(
        inst_data_MEM_data[117]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__21_ ( .D(n2504), .CLK(clk), .Q(
        inst_data_MEM_data[245]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__21_ ( .D(n2480), .CLK(clk), .Q(
        inst_data_MEM_data[213]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_21_ ( .D(inst_ID2EX_reg_N60), .CLK(
        clk), .Q(reg_read_data_1_EX[21]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_21_ ( .D(inst_EX2MEM_reg_N60), .CLK(
        clk), .Q(alu_result_MEM[21]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_21_ ( .D(u_MEM2WB_reg_N60), .CLK(clk), 
        .Q(alu_result_WB[21]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_22_ ( .D(u_MEM2WB_reg_N29), .CLK(clk), 
        .Q(mem_read_data_WB[22]) );
  DFFPOSX1 inst_register_registers_reg_7__22_ ( .D(n2447), .CLK(clk), .Q(
        inst_register_registers[246]) );
  DFFPOSX1 inst_register_registers_reg_6__22_ ( .D(n2423), .CLK(clk), .Q(
        inst_register_registers[214]) );
  DFFPOSX1 inst_register_registers_reg_5__22_ ( .D(n2384), .CLK(clk), .Q(
        inst_register_registers[182]) );
  DFFPOSX1 inst_register_registers_reg_4__22_ ( .D(n2352), .CLK(clk), .Q(
        inst_register_registers[150]) );
  DFFPOSX1 inst_register_registers_reg_3__22_ ( .D(n2323), .CLK(clk), .Q(
        inst_register_registers[118]) );
  DFFPOSX1 inst_register_registers_reg_2__22_ ( .D(n2287), .CLK(clk), .Q(
        inst_register_registers[86]) );
  DFFPOSX1 inst_register_registers_reg_1__22_ ( .D(n2255), .CLK(clk), .Q(
        inst_register_registers[54]) );
  DFFPOSX1 inst_register_registers_reg_0__22_ ( .D(n2223), .CLK(clk), .Q(
        inst_register_registers[22]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_22_ ( .D(inst_ID2EX_reg_N93), .CLK(
        clk), .Q(reg_read_data_2_EX[22]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_22_ ( .D(inst_EX2MEM_reg_N93), 
        .CLK(clk), .Q(write_mem_data_MEM[22]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__22_ ( .D(n2699), .CLK(clk), .Q(
        inst_data_MEM_data[86]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__22_ ( .D(n2667), .CLK(clk), .Q(
        inst_data_MEM_data[54]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__22_ ( .D(n2635), .CLK(clk), .Q(
        inst_data_MEM_data[22]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__22_ ( .D(n2596), .CLK(clk), .Q(
        inst_data_MEM_data[182]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__22_ ( .D(n2564), .CLK(clk), .Q(
        inst_data_MEM_data[150]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__22_ ( .D(n2535), .CLK(clk), .Q(
        inst_data_MEM_data[118]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__22_ ( .D(n2503), .CLK(clk), .Q(
        inst_data_MEM_data[246]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__22_ ( .D(n2479), .CLK(clk), .Q(
        inst_data_MEM_data[214]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_22_ ( .D(inst_ID2EX_reg_N61), .CLK(
        clk), .Q(reg_read_data_1_EX[22]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_22_ ( .D(inst_EX2MEM_reg_N61), .CLK(
        clk), .Q(alu_result_MEM[22]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_22_ ( .D(u_MEM2WB_reg_N61), .CLK(clk), 
        .Q(alu_result_WB[22]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_23_ ( .D(u_MEM2WB_reg_N30), .CLK(clk), 
        .Q(mem_read_data_WB[23]) );
  DFFPOSX1 inst_register_registers_reg_7__23_ ( .D(n2446), .CLK(clk), .Q(
        inst_register_registers[247]) );
  DFFPOSX1 inst_register_registers_reg_6__23_ ( .D(n2422), .CLK(clk), .Q(
        inst_register_registers[215]) );
  DFFPOSX1 inst_register_registers_reg_5__23_ ( .D(n2383), .CLK(clk), .Q(
        inst_register_registers[183]) );
  DFFPOSX1 inst_register_registers_reg_4__23_ ( .D(n2351), .CLK(clk), .Q(
        inst_register_registers[151]) );
  DFFPOSX1 inst_register_registers_reg_3__23_ ( .D(n2322), .CLK(clk), .Q(
        inst_register_registers[119]) );
  DFFPOSX1 inst_register_registers_reg_2__23_ ( .D(n2286), .CLK(clk), .Q(
        inst_register_registers[87]) );
  DFFPOSX1 inst_register_registers_reg_1__23_ ( .D(n2254), .CLK(clk), .Q(
        inst_register_registers[55]) );
  DFFPOSX1 inst_register_registers_reg_0__23_ ( .D(n2222), .CLK(clk), .Q(
        inst_register_registers[23]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_23_ ( .D(inst_ID2EX_reg_N94), .CLK(
        clk), .Q(reg_read_data_2_EX[23]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_23_ ( .D(inst_EX2MEM_reg_N94), 
        .CLK(clk), .Q(write_mem_data_MEM[23]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__23_ ( .D(n2698), .CLK(clk), .Q(
        inst_data_MEM_data[87]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__23_ ( .D(n2666), .CLK(clk), .Q(
        inst_data_MEM_data[55]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__23_ ( .D(n2634), .CLK(clk), .Q(
        inst_data_MEM_data[23]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__23_ ( .D(n2595), .CLK(clk), .Q(
        inst_data_MEM_data[183]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__23_ ( .D(n2563), .CLK(clk), .Q(
        inst_data_MEM_data[151]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__23_ ( .D(n2534), .CLK(clk), .Q(
        inst_data_MEM_data[119]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__23_ ( .D(n2502), .CLK(clk), .Q(
        inst_data_MEM_data[247]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__23_ ( .D(n2478), .CLK(clk), .Q(
        inst_data_MEM_data[215]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_23_ ( .D(inst_ID2EX_reg_N62), .CLK(
        clk), .Q(reg_read_data_1_EX[23]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_23_ ( .D(inst_EX2MEM_reg_N62), .CLK(
        clk), .Q(alu_result_MEM[23]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_23_ ( .D(u_MEM2WB_reg_N62), .CLK(clk), 
        .Q(alu_result_WB[23]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_24_ ( .D(u_MEM2WB_reg_N31), .CLK(clk), 
        .Q(mem_read_data_WB[24]) );
  DFFPOSX1 inst_register_registers_reg_7__24_ ( .D(n2445), .CLK(clk), .Q(
        inst_register_registers[248]) );
  DFFPOSX1 inst_register_registers_reg_6__24_ ( .D(n2421), .CLK(clk), .Q(
        inst_register_registers[216]) );
  DFFPOSX1 inst_register_registers_reg_5__24_ ( .D(n2382), .CLK(clk), .Q(
        inst_register_registers[184]) );
  DFFPOSX1 inst_register_registers_reg_4__24_ ( .D(n2350), .CLK(clk), .Q(
        inst_register_registers[152]) );
  DFFPOSX1 inst_register_registers_reg_3__24_ ( .D(n2321), .CLK(clk), .Q(
        inst_register_registers[120]) );
  DFFPOSX1 inst_register_registers_reg_2__24_ ( .D(n2285), .CLK(clk), .Q(
        inst_register_registers[88]) );
  DFFPOSX1 inst_register_registers_reg_1__24_ ( .D(n2253), .CLK(clk), .Q(
        inst_register_registers[56]) );
  DFFPOSX1 inst_register_registers_reg_0__24_ ( .D(n2221), .CLK(clk), .Q(
        inst_register_registers[24]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_24_ ( .D(inst_ID2EX_reg_N95), .CLK(
        clk), .Q(reg_read_data_2_EX[24]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_24_ ( .D(inst_EX2MEM_reg_N95), 
        .CLK(clk), .Q(write_mem_data_MEM[24]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__24_ ( .D(n2697), .CLK(clk), .Q(
        inst_data_MEM_data[88]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__24_ ( .D(n2665), .CLK(clk), .Q(
        inst_data_MEM_data[56]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__24_ ( .D(n2633), .CLK(clk), .Q(
        inst_data_MEM_data[24]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__24_ ( .D(n2594), .CLK(clk), .Q(
        inst_data_MEM_data[184]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__24_ ( .D(n2562), .CLK(clk), .Q(
        inst_data_MEM_data[152]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__24_ ( .D(n2533), .CLK(clk), .Q(
        inst_data_MEM_data[120]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__24_ ( .D(n2501), .CLK(clk), .Q(
        inst_data_MEM_data[248]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__24_ ( .D(n2477), .CLK(clk), .Q(
        inst_data_MEM_data[216]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_24_ ( .D(inst_ID2EX_reg_N63), .CLK(
        clk), .Q(reg_read_data_1_EX[24]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_24_ ( .D(inst_EX2MEM_reg_N63), .CLK(
        clk), .Q(alu_result_MEM[24]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_24_ ( .D(u_MEM2WB_reg_N63), .CLK(clk), 
        .Q(alu_result_WB[24]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_25_ ( .D(u_MEM2WB_reg_N32), .CLK(clk), 
        .Q(mem_read_data_WB[25]) );
  DFFPOSX1 inst_register_registers_reg_7__25_ ( .D(n2444), .CLK(clk), .Q(
        inst_register_registers[249]) );
  DFFPOSX1 inst_register_registers_reg_6__25_ ( .D(n2420), .CLK(clk), .Q(
        inst_register_registers[217]) );
  DFFPOSX1 inst_register_registers_reg_5__25_ ( .D(n2381), .CLK(clk), .Q(
        inst_register_registers[185]) );
  DFFPOSX1 inst_register_registers_reg_4__25_ ( .D(n2349), .CLK(clk), .Q(
        inst_register_registers[153]) );
  DFFPOSX1 inst_register_registers_reg_3__25_ ( .D(n2320), .CLK(clk), .Q(
        inst_register_registers[121]) );
  DFFPOSX1 inst_register_registers_reg_2__25_ ( .D(n2284), .CLK(clk), .Q(
        inst_register_registers[89]) );
  DFFPOSX1 inst_register_registers_reg_1__25_ ( .D(n2252), .CLK(clk), .Q(
        inst_register_registers[57]) );
  DFFPOSX1 inst_register_registers_reg_0__25_ ( .D(n2220), .CLK(clk), .Q(
        inst_register_registers[25]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_25_ ( .D(inst_ID2EX_reg_N96), .CLK(
        clk), .Q(reg_read_data_2_EX[25]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_25_ ( .D(inst_EX2MEM_reg_N96), 
        .CLK(clk), .Q(write_mem_data_MEM[25]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__25_ ( .D(n2696), .CLK(clk), .Q(
        inst_data_MEM_data[89]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__25_ ( .D(n2664), .CLK(clk), .Q(
        inst_data_MEM_data[57]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__25_ ( .D(n2632), .CLK(clk), .Q(
        inst_data_MEM_data[25]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__25_ ( .D(n2593), .CLK(clk), .Q(
        inst_data_MEM_data[185]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__25_ ( .D(n2561), .CLK(clk), .Q(
        inst_data_MEM_data[153]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__25_ ( .D(n2532), .CLK(clk), .Q(
        inst_data_MEM_data[121]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__25_ ( .D(n2500), .CLK(clk), .Q(
        inst_data_MEM_data[249]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__25_ ( .D(n2476), .CLK(clk), .Q(
        inst_data_MEM_data[217]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_25_ ( .D(inst_ID2EX_reg_N64), .CLK(
        clk), .Q(reg_read_data_1_EX[25]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_25_ ( .D(inst_EX2MEM_reg_N64), .CLK(
        clk), .Q(alu_result_MEM[25]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_25_ ( .D(u_MEM2WB_reg_N64), .CLK(clk), 
        .Q(alu_result_WB[25]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_26_ ( .D(u_MEM2WB_reg_N33), .CLK(clk), 
        .Q(mem_read_data_WB[26]) );
  DFFPOSX1 inst_register_registers_reg_7__26_ ( .D(n2443), .CLK(clk), .Q(
        inst_register_registers[250]) );
  DFFPOSX1 inst_register_registers_reg_6__26_ ( .D(n2419), .CLK(clk), .Q(
        inst_register_registers[218]) );
  DFFPOSX1 inst_register_registers_reg_5__26_ ( .D(n2380), .CLK(clk), .Q(
        inst_register_registers[186]) );
  DFFPOSX1 inst_register_registers_reg_4__26_ ( .D(n2348), .CLK(clk), .Q(
        inst_register_registers[154]) );
  DFFPOSX1 inst_register_registers_reg_3__26_ ( .D(n2319), .CLK(clk), .Q(
        inst_register_registers[122]) );
  DFFPOSX1 inst_register_registers_reg_2__26_ ( .D(n2283), .CLK(clk), .Q(
        inst_register_registers[90]) );
  DFFPOSX1 inst_register_registers_reg_1__26_ ( .D(n2251), .CLK(clk), .Q(
        inst_register_registers[58]) );
  DFFPOSX1 inst_register_registers_reg_0__26_ ( .D(n2219), .CLK(clk), .Q(
        inst_register_registers[26]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_26_ ( .D(inst_ID2EX_reg_N97), .CLK(
        clk), .Q(reg_read_data_2_EX[26]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_26_ ( .D(inst_EX2MEM_reg_N97), 
        .CLK(clk), .Q(write_mem_data_MEM[26]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__26_ ( .D(n2695), .CLK(clk), .Q(
        inst_data_MEM_data[90]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__26_ ( .D(n2663), .CLK(clk), .Q(
        inst_data_MEM_data[58]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__26_ ( .D(n2631), .CLK(clk), .Q(
        inst_data_MEM_data[26]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__26_ ( .D(n2592), .CLK(clk), .Q(
        inst_data_MEM_data[186]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__26_ ( .D(n2560), .CLK(clk), .Q(
        inst_data_MEM_data[154]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__26_ ( .D(n2531), .CLK(clk), .Q(
        inst_data_MEM_data[122]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__26_ ( .D(n2499), .CLK(clk), .Q(
        inst_data_MEM_data[250]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__26_ ( .D(n2475), .CLK(clk), .Q(
        inst_data_MEM_data[218]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_26_ ( .D(inst_ID2EX_reg_N65), .CLK(
        clk), .Q(reg_read_data_1_EX[26]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_26_ ( .D(inst_EX2MEM_reg_N65), .CLK(
        clk), .Q(alu_result_MEM[26]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_26_ ( .D(u_MEM2WB_reg_N65), .CLK(clk), 
        .Q(alu_result_WB[26]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_27_ ( .D(u_MEM2WB_reg_N34), .CLK(clk), 
        .Q(mem_read_data_WB[27]) );
  DFFPOSX1 inst_register_registers_reg_7__27_ ( .D(n2442), .CLK(clk), .Q(
        inst_register_registers[251]) );
  DFFPOSX1 inst_register_registers_reg_6__27_ ( .D(n2418), .CLK(clk), .Q(
        inst_register_registers[219]) );
  DFFPOSX1 inst_register_registers_reg_5__27_ ( .D(n2379), .CLK(clk), .Q(
        inst_register_registers[187]) );
  DFFPOSX1 inst_register_registers_reg_4__27_ ( .D(n2347), .CLK(clk), .Q(
        inst_register_registers[155]) );
  DFFPOSX1 inst_register_registers_reg_3__27_ ( .D(n2318), .CLK(clk), .Q(
        inst_register_registers[123]) );
  DFFPOSX1 inst_register_registers_reg_2__27_ ( .D(n2282), .CLK(clk), .Q(
        inst_register_registers[91]) );
  DFFPOSX1 inst_register_registers_reg_1__27_ ( .D(n2250), .CLK(clk), .Q(
        inst_register_registers[59]) );
  DFFPOSX1 inst_register_registers_reg_0__27_ ( .D(n2218), .CLK(clk), .Q(
        inst_register_registers[27]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_27_ ( .D(inst_ID2EX_reg_N98), .CLK(
        clk), .Q(reg_read_data_2_EX[27]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_27_ ( .D(inst_EX2MEM_reg_N98), 
        .CLK(clk), .Q(write_mem_data_MEM[27]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__27_ ( .D(n2694), .CLK(clk), .Q(
        inst_data_MEM_data[91]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__27_ ( .D(n2662), .CLK(clk), .Q(
        inst_data_MEM_data[59]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__27_ ( .D(n2630), .CLK(clk), .Q(
        inst_data_MEM_data[27]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__27_ ( .D(n2591), .CLK(clk), .Q(
        inst_data_MEM_data[187]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__27_ ( .D(n2559), .CLK(clk), .Q(
        inst_data_MEM_data[155]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__27_ ( .D(n2530), .CLK(clk), .Q(
        inst_data_MEM_data[123]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__27_ ( .D(n2498), .CLK(clk), .Q(
        inst_data_MEM_data[251]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__27_ ( .D(n2474), .CLK(clk), .Q(
        inst_data_MEM_data[219]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_27_ ( .D(inst_ID2EX_reg_N66), .CLK(
        clk), .Q(reg_read_data_1_EX[27]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_27_ ( .D(inst_EX2MEM_reg_N66), .CLK(
        clk), .Q(alu_result_MEM[27]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_27_ ( .D(u_MEM2WB_reg_N66), .CLK(clk), 
        .Q(alu_result_WB[27]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_28_ ( .D(u_MEM2WB_reg_N35), .CLK(clk), 
        .Q(mem_read_data_WB[28]) );
  DFFPOSX1 inst_register_registers_reg_7__28_ ( .D(n2441), .CLK(clk), .Q(
        inst_register_registers[252]) );
  DFFPOSX1 inst_register_registers_reg_6__28_ ( .D(n2417), .CLK(clk), .Q(
        inst_register_registers[220]) );
  DFFPOSX1 inst_register_registers_reg_5__28_ ( .D(n2378), .CLK(clk), .Q(
        inst_register_registers[188]) );
  DFFPOSX1 inst_register_registers_reg_4__28_ ( .D(n2346), .CLK(clk), .Q(
        inst_register_registers[156]) );
  DFFPOSX1 inst_register_registers_reg_3__28_ ( .D(n2317), .CLK(clk), .Q(
        inst_register_registers[124]) );
  DFFPOSX1 inst_register_registers_reg_2__28_ ( .D(n2281), .CLK(clk), .Q(
        inst_register_registers[92]) );
  DFFPOSX1 inst_register_registers_reg_1__28_ ( .D(n2249), .CLK(clk), .Q(
        inst_register_registers[60]) );
  DFFPOSX1 inst_register_registers_reg_0__28_ ( .D(n2217), .CLK(clk), .Q(
        inst_register_registers[28]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_28_ ( .D(inst_ID2EX_reg_N99), .CLK(
        clk), .Q(reg_read_data_2_EX[28]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_28_ ( .D(inst_EX2MEM_reg_N99), 
        .CLK(clk), .Q(write_mem_data_MEM[28]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__28_ ( .D(n2693), .CLK(clk), .Q(
        inst_data_MEM_data[92]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__28_ ( .D(n2661), .CLK(clk), .Q(
        inst_data_MEM_data[60]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__28_ ( .D(n2629), .CLK(clk), .Q(
        inst_data_MEM_data[28]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__28_ ( .D(n2590), .CLK(clk), .Q(
        inst_data_MEM_data[188]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__28_ ( .D(n2558), .CLK(clk), .Q(
        inst_data_MEM_data[156]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__28_ ( .D(n2529), .CLK(clk), .Q(
        inst_data_MEM_data[124]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__28_ ( .D(n2497), .CLK(clk), .Q(
        inst_data_MEM_data[252]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__28_ ( .D(n2473), .CLK(clk), .Q(
        inst_data_MEM_data[220]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_28_ ( .D(inst_ID2EX_reg_N67), .CLK(
        clk), .Q(reg_read_data_1_EX[28]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_28_ ( .D(inst_EX2MEM_reg_N67), .CLK(
        clk), .Q(alu_result_MEM[28]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_28_ ( .D(u_MEM2WB_reg_N67), .CLK(clk), 
        .Q(alu_result_WB[28]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_29_ ( .D(u_MEM2WB_reg_N36), .CLK(clk), 
        .Q(mem_read_data_WB[29]) );
  DFFPOSX1 inst_register_registers_reg_7__29_ ( .D(n2470), .CLK(clk), .Q(
        inst_register_registers[253]) );
  DFFPOSX1 inst_register_registers_reg_6__29_ ( .D(n2416), .CLK(clk), .Q(
        inst_register_registers[221]) );
  DFFPOSX1 inst_register_registers_reg_5__29_ ( .D(n2377), .CLK(clk), .Q(
        inst_register_registers[189]) );
  DFFPOSX1 inst_register_registers_reg_4__29_ ( .D(n2345), .CLK(clk), .Q(
        inst_register_registers[157]) );
  DFFPOSX1 inst_register_registers_reg_3__29_ ( .D(n2316), .CLK(clk), .Q(
        inst_register_registers[125]) );
  DFFPOSX1 inst_register_registers_reg_2__29_ ( .D(n2280), .CLK(clk), .Q(
        inst_register_registers[93]) );
  DFFPOSX1 inst_register_registers_reg_1__29_ ( .D(n2248), .CLK(clk), .Q(
        inst_register_registers[61]) );
  DFFPOSX1 inst_register_registers_reg_0__29_ ( .D(n2216), .CLK(clk), .Q(
        inst_register_registers[29]) );
  DFFPOSX1 inst_ID2EX_reg_register_2_reg_29_ ( .D(inst_ID2EX_reg_N100), .CLK(
        clk), .Q(reg_read_data_2_EX[29]) );
  DFFPOSX1 inst_EX2MEM_reg_write_mem_data_reg_29_ ( .D(inst_EX2MEM_reg_N100), 
        .CLK(clk), .Q(write_mem_data_MEM[29]) );
  DFFPOSX1 inst_data_MEM_data_reg_2__29_ ( .D(n2692), .CLK(clk), .Q(
        inst_data_MEM_data[93]) );
  DFFPOSX1 inst_data_MEM_data_reg_1__29_ ( .D(n2660), .CLK(clk), .Q(
        inst_data_MEM_data[61]) );
  DFFPOSX1 inst_data_MEM_data_reg_0__29_ ( .D(n2628), .CLK(clk), .Q(
        inst_data_MEM_data[29]) );
  DFFPOSX1 inst_data_MEM_data_reg_5__29_ ( .D(n2589), .CLK(clk), .Q(
        inst_data_MEM_data[189]) );
  DFFPOSX1 inst_data_MEM_data_reg_4__29_ ( .D(n2557), .CLK(clk), .Q(
        inst_data_MEM_data[157]) );
  DFFPOSX1 inst_data_MEM_data_reg_3__29_ ( .D(n2528), .CLK(clk), .Q(
        inst_data_MEM_data[125]) );
  DFFPOSX1 inst_data_MEM_data_reg_7__29_ ( .D(n2526), .CLK(clk), .Q(
        inst_data_MEM_data[253]) );
  DFFPOSX1 inst_data_MEM_data_reg_6__29_ ( .D(n2472), .CLK(clk), .Q(
        inst_data_MEM_data[221]) );
  DFFPOSX1 inst_ID2EX_reg_register_1_reg_29_ ( .D(inst_ID2EX_reg_N68), .CLK(
        clk), .Q(reg_read_data_1_EX[29]) );
  DFFPOSX1 inst_EX2MEM_reg_alu_result_reg_29_ ( .D(inst_EX2MEM_reg_N68), .CLK(
        clk), .Q(alu_result_MEM[29]) );
  DFFPOSX1 u_MEM2WB_reg_alu_result_reg_29_ ( .D(u_MEM2WB_reg_N68), .CLK(clk), 
        .Q(alu_result_WB[29]) );
  DFFPOSX1 u_MEM2WB_reg_read_data_reg_30_ ( .D(u_MEM2WB_reg_N37), .CLK(clk), 
        .Q(mem_read_data_WB[30]) );
  DFFPOSX1 inst_PC_inst_addr_reg_0_ ( .D(n2214), .CLK(clk), .Q(inst_address[0]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_0_ ( .D(n2727), .CLK(clk), .Q(
        inst_addr_ID[0]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_0_ ( .D(inst_ID2EX_reg_N7), .CLK(clk), 
        .Q(shifted_address_EX[0]) );
  DFFPOSX1 inst_PC_inst_addr_reg_1_ ( .D(n2213), .CLK(clk), .Q(inst_address[1]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_1_ ( .D(n2728), .CLK(clk), .Q(
        inst_addr_ID[1]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_1_ ( .D(inst_ID2EX_reg_N8), .CLK(clk), 
        .Q(shifted_address_EX[1]) );
  DFFPOSX1 inst_PC_inst_addr_reg_2_ ( .D(n2212), .CLK(clk), .Q(inst_address[2]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_2_ ( .D(n2729), .CLK(clk), .Q(
        inst_addr_ID[2]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_2_ ( .D(inst_ID2EX_reg_N9), .CLK(clk), 
        .Q(inst_addr_EX[2]) );
  DFFPOSX1 inst_PC_inst_addr_reg_3_ ( .D(n2211), .CLK(clk), .Q(inst_address[3]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_3_ ( .D(n2730), .CLK(clk), .Q(
        inst_addr_ID[3]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_3_ ( .D(inst_ID2EX_reg_N10), .CLK(clk), 
        .Q(inst_addr_EX[3]) );
  DFFPOSX1 inst_PC_inst_addr_reg_4_ ( .D(n2210), .CLK(clk), .Q(inst_address[4]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_4_ ( .D(n2731), .CLK(clk), .Q(
        inst_addr_ID[4]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_4_ ( .D(inst_ID2EX_reg_N11), .CLK(clk), 
        .Q(inst_addr_EX[4]) );
  DFFPOSX1 inst_PC_inst_addr_reg_5_ ( .D(n2209), .CLK(clk), .Q(inst_address[5]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_5_ ( .D(n2732), .CLK(clk), .Q(
        inst_addr_ID[5]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_5_ ( .D(inst_ID2EX_reg_N12), .CLK(clk), 
        .Q(inst_addr_EX[5]) );
  DFFPOSX1 inst_PC_inst_addr_reg_6_ ( .D(n2208), .CLK(clk), .Q(inst_address[6]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_6_ ( .D(n2733), .CLK(clk), .Q(
        inst_addr_ID[6]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_6_ ( .D(inst_ID2EX_reg_N13), .CLK(clk), 
        .Q(inst_addr_EX[6]) );
  DFFPOSX1 inst_PC_inst_addr_reg_7_ ( .D(n2207), .CLK(clk), .Q(inst_address[7]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_7_ ( .D(n2734), .CLK(clk), .Q(
        inst_addr_ID[7]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_7_ ( .D(inst_ID2EX_reg_N14), .CLK(clk), 
        .Q(inst_addr_EX[7]) );
  DFFPOSX1 inst_PC_inst_addr_reg_8_ ( .D(n2206), .CLK(clk), .Q(inst_address[8]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_8_ ( .D(n2735), .CLK(clk), .Q(
        inst_addr_ID[8]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_8_ ( .D(inst_ID2EX_reg_N15), .CLK(clk), 
        .Q(inst_addr_EX[8]) );
  DFFPOSX1 inst_PC_inst_addr_reg_9_ ( .D(n2205), .CLK(clk), .Q(inst_address[9]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_9_ ( .D(n2736), .CLK(clk), .Q(
        inst_addr_ID[9]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_9_ ( .D(inst_ID2EX_reg_N16), .CLK(clk), 
        .Q(inst_addr_EX[9]) );
  DFFPOSX1 inst_PC_inst_addr_reg_10_ ( .D(n2204), .CLK(clk), .Q(
        inst_address[10]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_10_ ( .D(n2737), .CLK(clk), .Q(
        inst_addr_ID[10]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_10_ ( .D(inst_ID2EX_reg_N17), .CLK(clk), 
        .Q(inst_addr_EX[10]) );
  DFFPOSX1 inst_PC_inst_addr_reg_11_ ( .D(n2203), .CLK(clk), .Q(
        inst_address[11]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_11_ ( .D(n2738), .CLK(clk), .Q(
        inst_addr_ID[11]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_11_ ( .D(inst_ID2EX_reg_N18), .CLK(clk), 
        .Q(inst_addr_EX[11]) );
  DFFPOSX1 inst_PC_inst_addr_reg_12_ ( .D(n2202), .CLK(clk), .Q(
        inst_address[12]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_12_ ( .D(n2739), .CLK(clk), .Q(
        inst_addr_ID[12]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_12_ ( .D(inst_ID2EX_reg_N19), .CLK(clk), 
        .Q(inst_addr_EX[12]) );
  DFFPOSX1 inst_PC_inst_addr_reg_13_ ( .D(n2201), .CLK(clk), .Q(
        inst_address[13]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_13_ ( .D(n2740), .CLK(clk), .Q(
        inst_addr_ID[13]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_13_ ( .D(inst_ID2EX_reg_N20), .CLK(clk), 
        .Q(inst_addr_EX[13]) );
  DFFPOSX1 inst_PC_inst_addr_reg_14_ ( .D(n2200), .CLK(clk), .Q(
        inst_address[14]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_14_ ( .D(n2741), .CLK(clk), .Q(
        inst_addr_ID[14]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_14_ ( .D(inst_ID2EX_reg_N21), .CLK(clk), 
        .Q(inst_addr_EX[14]) );
  DFFPOSX1 inst_PC_inst_addr_reg_15_ ( .D(n2199), .CLK(clk), .Q(
        inst_address[15]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_15_ ( .D(n2742), .CLK(clk), .Q(
        inst_addr_ID[15]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_15_ ( .D(inst_ID2EX_reg_N22), .CLK(clk), 
        .Q(inst_addr_EX[15]) );
  DFFPOSX1 inst_PC_inst_addr_reg_16_ ( .D(n2198), .CLK(clk), .Q(
        inst_address[16]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_16_ ( .D(n2743), .CLK(clk), .Q(
        inst_addr_ID[16]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_16_ ( .D(inst_ID2EX_reg_N23), .CLK(clk), 
        .Q(inst_addr_EX[16]) );
  DFFPOSX1 inst_PC_inst_addr_reg_17_ ( .D(n2197), .CLK(clk), .Q(
        inst_address[17]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_17_ ( .D(n2744), .CLK(clk), .Q(
        inst_addr_ID[17]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_17_ ( .D(inst_ID2EX_reg_N24), .CLK(clk), 
        .Q(inst_addr_EX[17]) );
  DFFPOSX1 inst_PC_inst_addr_reg_18_ ( .D(n2196), .CLK(clk), .Q(
        inst_address[18]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_18_ ( .D(n2745), .CLK(clk), .Q(
        inst_addr_ID[18]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_18_ ( .D(inst_ID2EX_reg_N25), .CLK(clk), 
        .Q(inst_addr_EX[18]) );
  DFFPOSX1 inst_PC_inst_addr_reg_19_ ( .D(n2195), .CLK(clk), .Q(
        inst_address[19]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_19_ ( .D(n2746), .CLK(clk), .Q(
        inst_addr_ID[19]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_19_ ( .D(inst_ID2EX_reg_N26), .CLK(clk), 
        .Q(inst_addr_EX[19]) );
  DFFPOSX1 inst_PC_inst_addr_reg_20_ ( .D(n2194), .CLK(clk), .Q(
        inst_address[20]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_20_ ( .D(n2747), .CLK(clk), .Q(
        inst_addr_ID[20]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_20_ ( .D(inst_ID2EX_reg_N27), .CLK(clk), 
        .Q(inst_addr_EX[20]) );
  DFFPOSX1 inst_PC_inst_addr_reg_21_ ( .D(n2193), .CLK(clk), .Q(
        inst_address[21]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_21_ ( .D(n2748), .CLK(clk), .Q(
        inst_addr_ID[21]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_21_ ( .D(inst_ID2EX_reg_N28), .CLK(clk), 
        .Q(inst_addr_EX[21]) );
  DFFPOSX1 inst_PC_inst_addr_reg_22_ ( .D(n2192), .CLK(clk), .Q(
        inst_address[22]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_22_ ( .D(n2749), .CLK(clk), .Q(
        inst_addr_ID[22]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_22_ ( .D(inst_ID2EX_reg_N29), .CLK(clk), 
        .Q(inst_addr_EX[22]) );
  DFFPOSX1 inst_PC_inst_addr_reg_23_ ( .D(n2191), .CLK(clk), .Q(
        inst_address[23]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_23_ ( .D(n2750), .CLK(clk), .Q(
        inst_addr_ID[23]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_23_ ( .D(inst_ID2EX_reg_N30), .CLK(clk), 
        .Q(inst_addr_EX[23]) );
  DFFPOSX1 inst_PC_inst_addr_reg_24_ ( .D(n2190), .CLK(clk), .Q(
        inst_address[24]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_24_ ( .D(n2751), .CLK(clk), .Q(
        inst_addr_ID[24]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_24_ ( .D(inst_ID2EX_reg_N31), .CLK(clk), 
        .Q(inst_addr_EX[24]) );
  DFFPOSX1 inst_PC_inst_addr_reg_25_ ( .D(n2189), .CLK(clk), .Q(
        inst_address[25]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_25_ ( .D(n2752), .CLK(clk), .Q(
        inst_addr_ID[25]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_25_ ( .D(inst_ID2EX_reg_N32), .CLK(clk), 
        .Q(inst_addr_EX[25]) );
  DFFPOSX1 inst_PC_inst_addr_reg_26_ ( .D(n2188), .CLK(clk), .Q(
        inst_address[26]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_26_ ( .D(n2753), .CLK(clk), .Q(
        inst_addr_ID[26]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_26_ ( .D(inst_ID2EX_reg_N33), .CLK(clk), 
        .Q(inst_addr_EX[26]) );
  DFFPOSX1 inst_PC_inst_addr_reg_27_ ( .D(n2187), .CLK(clk), .Q(
        inst_address[27]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_27_ ( .D(n2754), .CLK(clk), .Q(
        inst_addr_ID[27]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_27_ ( .D(inst_ID2EX_reg_N34), .CLK(clk), 
        .Q(inst_addr_EX[27]) );
  DFFPOSX1 inst_PC_inst_addr_reg_28_ ( .D(n2186), .CLK(clk), .Q(
        inst_address[28]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_28_ ( .D(n2755), .CLK(clk), .Q(
        inst_addr_ID[28]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_28_ ( .D(inst_ID2EX_reg_N35), .CLK(clk), 
        .Q(inst_addr_EX[28]) );
  DFFPOSX1 inst_PC_inst_addr_reg_29_ ( .D(n2185), .CLK(clk), .Q(
        inst_address[29]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_29_ ( .D(n2756), .CLK(clk), .Q(
        inst_addr_ID[29]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_29_ ( .D(inst_ID2EX_reg_N36), .CLK(clk), 
        .Q(inst_addr_EX[29]) );
  DFFPOSX1 inst_PC_inst_addr_reg_30_ ( .D(n2183), .CLK(clk), .Q(
        inst_address[30]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_30_ ( .D(n2757), .CLK(clk), .Q(
        inst_addr_ID[30]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_30_ ( .D(inst_ID2EX_reg_N37), .CLK(clk), 
        .Q(inst_addr_EX[30]) );
  DFFPOSX1 inst_PC_inst_addr_reg_31_ ( .D(n2791), .CLK(clk), .Q(
        inst_address[31]) );
  DFFPOSX1 inst_IF2ID_reg_inst_address_reg_31_ ( .D(n2758), .CLK(clk), .Q(
        inst_addr_ID[31]) );
  DFFPOSX1 inst_ID2EX_reg_address_reg_31_ ( .D(inst_ID2EX_reg_N38), .CLK(clk), 
        .Q(inst_addr_EX[31]) );
  INVX4 U3191 ( .A(n4050), .Y(n4263) );
  INVX1 U3192 ( .A(n4171), .Y(n4152) );
  INVX1 U3193 ( .A(n4150), .Y(n4206) );
  INVX1 U3194 ( .A(n4189), .Y(n4163) );
  INVX1 U3195 ( .A(n3963), .Y(n4177) );
  AND2X2 U3196 ( .A(n3943), .B(n3727), .Y(n3728) );
  INVX1 U3197 ( .A(n5198), .Y(n5199) );
  INVX1 U3198 ( .A(n5195), .Y(n5196) );
  INVX1 U3199 ( .A(n4968), .Y(n4931) );
  INVX1 U3200 ( .A(n4925), .Y(n4889) );
  INVX1 U3201 ( .A(n4832), .Y(n4796) );
  INVX1 U3202 ( .A(shifted_address_MEM[17]), .Y(n4304) );
  INVX1 U3203 ( .A(shifted_address_MEM[3]), .Y(n4272) );
  BUFX2 U3204 ( .A(n4033), .Y(n4050) );
  INVX4 U3205 ( .A(n3933), .Y(n2795) );
  INVX4 U3206 ( .A(n4617), .Y(n4727) );
  BUFX2 U3207 ( .A(n4526), .Y(n4451) );
  BUFX2 U3208 ( .A(n4602), .Y(n4435) );
  BUFX2 U3209 ( .A(n4609), .Y(n4442) );
  BUFX2 U3210 ( .A(n4603), .Y(n4437) );
  INVX4 U3211 ( .A(n4705), .Y(n2796) );
  INVX1 U3212 ( .A(n4190), .Y(n4162) );
  INVX4 U3213 ( .A(n4515), .Y(n2797) );
  INVX4 U3214 ( .A(n4457), .Y(n2798) );
  INVX4 U3215 ( .A(n4474), .Y(n2799) );
  INVX4 U3216 ( .A(n4468), .Y(n2800) );
  AND2X2 U3217 ( .A(n3943), .B(n3730), .Y(n3731) );
  AND2X1 U3218 ( .A(n3943), .B(n3724), .Y(n3725) );
  BUFX2 U3219 ( .A(n3552), .Y(n3156) );
  BUFX2 U3220 ( .A(n3324), .Y(n3073) );
  BUFX2 U3221 ( .A(n3564), .Y(n3031) );
  BUFX2 U3222 ( .A(n3535), .Y(n3207) );
  BUFX2 U3223 ( .A(n3419), .Y(n3038) );
  BUFX2 U3224 ( .A(n3562), .Y(n3041) );
  BUFX2 U3225 ( .A(n3563), .Y(n3032) );
  BUFX2 U3226 ( .A(n3559), .Y(n3071) );
  INVX4 U3227 ( .A(n3223), .Y(n2801) );
  INVX4 U3228 ( .A(n3205), .Y(n2802) );
  INVX4 U3229 ( .A(n3208), .Y(n2803) );
  INVX4 U3230 ( .A(n3209), .Y(n2804) );
  INVX4 U3231 ( .A(n3381), .Y(n2805) );
  INVX4 U3232 ( .A(n3070), .Y(n2806) );
  INVX4 U3233 ( .A(n3245), .Y(n2807) );
  INVX4 U3234 ( .A(n3080), .Y(n2808) );
  INVX4 U3235 ( .A(n4426), .Y(n2809) );
  BUFX2 U3236 ( .A(n3733), .Y(n2901) );
  BUFX2 U3237 ( .A(n3537), .Y(n3148) );
  BUFX2 U3238 ( .A(n3561), .Y(n3030) );
  BUFX2 U3239 ( .A(n5345), .Y(n5317) );
  BUFX2 U3240 ( .A(n5386), .Y(n5355) );
  INVX4 U3241 ( .A(n5209), .Y(n2810) );
  INVX4 U3242 ( .A(n5155), .Y(n2811) );
  INVX4 U3243 ( .A(n5282), .Y(n2812) );
  INVX4 U3244 ( .A(n5437), .Y(n2813) );
  BUFX2 U3245 ( .A(n4870), .Y(n4836) );
  BUFX2 U3246 ( .A(n5486), .Y(n5430) );
  BUFX2 U3247 ( .A(n4966), .Y(n4929) );
  BUFX2 U3248 ( .A(n4923), .Y(n4887) );
  INVX4 U3249 ( .A(n5393), .Y(n5427) );
  INVX4 U3250 ( .A(n5244), .Y(n5278) );
  BUFX2 U3251 ( .A(n5313), .Y(n5280) );
  BUFX2 U3252 ( .A(n5388), .Y(n5354) );
  BUFX2 U3253 ( .A(n5351), .Y(n5316) );
  BUFX2 U3254 ( .A(n5240), .Y(n5203) );
  BUFX2 U3255 ( .A(n5234), .Y(n5120) );
  BUFX2 U3256 ( .A(n4830), .Y(n4797) );
  INVX2 U3257 ( .A(n5121), .Y(n5122) );
  INVX2 U3258 ( .A(n3949), .Y(n5204) );
  INVX4 U3259 ( .A(n2868), .Y(n2814) );
  INVX2 U3260 ( .A(n4872), .Y(n4835) );
  BUFX2 U3261 ( .A(n4792), .Y(n4760) );
  BUFX2 U3262 ( .A(n5000), .Y(n4754) );
  BUFX2 U3263 ( .A(n5112), .Y(n4878) );
  INVX1 U3264 ( .A(inst_address[6]), .Y(n4736) );
  INVX1 U3265 ( .A(inst_address[0]), .Y(n4747) );
  INVX1 U3266 ( .A(inst_address[1]), .Y(n4745) );
  INVX2 U3267 ( .A(n5392), .Y(n2815) );
  INVX2 U3268 ( .A(n3946), .Y(n3736) );
  INVX1 U3269 ( .A(n2924), .Y(n2925) );
  INVX1 U3270 ( .A(n2932), .Y(n2934) );
  OR2X1 U3271 ( .A(n3153), .B(n3154), .Y(n3245) );
  OR2X1 U3272 ( .A(n3153), .B(n3152), .Y(n3381) );
  OR2X1 U3273 ( .A(n3153), .B(n3151), .Y(n3208) );
  OR2X1 U3274 ( .A(n3151), .B(n3155), .Y(n3209) );
  OR2X1 U3275 ( .A(n3153), .B(n3149), .Y(n3205) );
  OR2X1 U3276 ( .A(n3155), .B(n3149), .Y(n3223) );
  OR2X1 U3277 ( .A(n3040), .B(n3034), .Y(n3070) );
  OR2X1 U3278 ( .A(n3035), .B(n3034), .Y(n3080) );
  INVX1 U3279 ( .A(n3852), .Y(n3847) );
  INVX1 U3280 ( .A(n3846), .Y(n3633) );
  INVX1 U3281 ( .A(n3854), .Y(n3632) );
  INVX1 U3282 ( .A(n3670), .Y(n5180) );
  INVX1 U3283 ( .A(n3674), .Y(n5178) );
  INVX1 U3284 ( .A(n3656), .Y(n5174) );
  INVX1 U3285 ( .A(n3389), .Y(n5167) );
  INVX1 U3286 ( .A(n3411), .Y(n5147) );
  OR2X1 U3287 ( .A(op_type_EX[2]), .B(n2838), .Y(n2839) );
  INVX1 U3288 ( .A(n4875), .Y(n4876) );
  INVX1 U3289 ( .A(n4757), .Y(n4758) );
  OR2X1 U3290 ( .A(n4445), .B(n4926), .Y(n4457) );
  INVX1 U3291 ( .A(n4750), .Y(n4751) );
  OR2X1 U3292 ( .A(n4445), .B(n4433), .Y(n4515) );
  INVX1 U3293 ( .A(n3594), .Y(n4927) );
  INVX1 U3294 ( .A(n3063), .Y(n3046) );
  OR2X1 U3295 ( .A(n2814), .B(n2869), .Y(n2870) );
  OR2X1 U3296 ( .A(n2896), .B(n2897), .Y(n2894) );
  OR2X1 U3297 ( .A(op_type_WB[3]), .B(n2843), .Y(n2844) );
  OR2X1 U3298 ( .A(n4445), .B(n4750), .Y(n4474) );
  OR2X1 U3299 ( .A(n4445), .B(n4875), .Y(n4468) );
  INVX1 U3300 ( .A(n5526), .Y(n4305) );
  INVX1 U3301 ( .A(n4139), .Y(n4056) );
  INVX1 U3302 ( .A(n2912), .Y(n2913) );
  INVX1 U3303 ( .A(n2916), .Y(n2917) );
  INVX1 U3304 ( .A(n2920), .Y(n2921) );
  INVX1 U3305 ( .A(n2937), .Y(n2938) );
  INVX1 U3306 ( .A(n2941), .Y(n2942) );
  INVX1 U3307 ( .A(n4926), .Y(n4928) );
  INVX1 U3308 ( .A(n4885), .Y(n4886) );
  INVX1 U3309 ( .A(n4833), .Y(n4834) );
  OR2X1 U3310 ( .A(n5392), .B(n3596), .Y(n5014) );
  INVX1 U3311 ( .A(n5061), .Y(n5009) );
  INVX1 U3312 ( .A(n3953), .Y(n4260) );
  INVX1 U3313 ( .A(n2969), .Y(n2970) );
  INVX1 U3314 ( .A(inst_addr_EX[29]), .Y(n4420) );
  INVX1 U3315 ( .A(inst_addr_EX[19]), .Y(n3628) );
  INVX1 U3316 ( .A(n5508), .Y(n5506) );
  OR2X1 U3317 ( .A(n3851), .B(n3639), .Y(n2200) );
  INVX1 U3318 ( .A(n4289), .Y(n3907) );
  INVX1 U3319 ( .A(n3543), .Y(inst_ID2EX_reg_N100) );
  INVX1 U3320 ( .A(n3337), .Y(inst_ID2EX_reg_N66) );
  INVX1 U3321 ( .A(n3237), .Y(inst_ID2EX_reg_N64) );
  INVX1 U3322 ( .A(n3222), .Y(inst_ID2EX_reg_N62) );
  INVX1 U3323 ( .A(n3215), .Y(inst_ID2EX_reg_N93) );
  INVX1 U3324 ( .A(n3244), .Y(inst_ID2EX_reg_N91) );
  INVX1 U3325 ( .A(n3504), .Y(inst_ID2EX_reg_N89) );
  INVX1 U3326 ( .A(n3351), .Y(inst_ID2EX_reg_N55) );
  INVX1 U3327 ( .A(n3512), .Y(inst_ID2EX_reg_N87) );
  INVX1 U3328 ( .A(n3365), .Y(inst_ID2EX_reg_N54) );
  INVX1 U3329 ( .A(n2985), .Y(inst_EX2MEM_reg_N53) );
  INVX1 U3330 ( .A(n3448), .Y(inst_ID2EX_reg_N85) );
  INVX1 U3331 ( .A(n3294), .Y(inst_ID2EX_reg_N52) );
  INVX1 U3332 ( .A(n2999), .Y(inst_EX2MEM_reg_N51) );
  INVX1 U3333 ( .A(n3136), .Y(inst_ID2EX_reg_N51) );
  INVX1 U3334 ( .A(n3020), .Y(inst_EX2MEM_reg_N49) );
  INVX1 U3335 ( .A(n3176), .Y(inst_ID2EX_reg_N49) );
  INVX1 U3336 ( .A(n3101), .Y(inst_ID2EX_reg_N48) );
  INVX1 U3337 ( .A(n3591), .Y(inst_EX2MEM_reg_N47) );
  INVX1 U3338 ( .A(n3069), .Y(inst_ID2EX_reg_N47) );
  INVX1 U3339 ( .A(n3122), .Y(inst_ID2EX_reg_N46) );
  INVX1 U3340 ( .A(n3432), .Y(inst_ID2EX_reg_N78) );
  INVX1 U3341 ( .A(n3129), .Y(inst_ID2EX_reg_N45) );
  INVX1 U3342 ( .A(n3402), .Y(inst_ID2EX_reg_N76) );
  INVX1 U3343 ( .A(n3190), .Y(inst_ID2EX_reg_N43) );
  INVX1 U3344 ( .A(n3183), .Y(inst_ID2EX_reg_N42) );
  INVX1 U3345 ( .A(n3597), .Y(n2522) );
  INVX1 U3346 ( .A(n3490), .Y(inst_ID2EX_reg_N74) );
  INVX1 U3347 ( .A(n4044), .Y(n4051) );
  INVX1 U3348 ( .A(n3519), .Y(inst_ID2EX_reg_N72) );
  INVX1 U3349 ( .A(n4036), .Y(n4041) );
  INVX1 U3350 ( .A(n3455), .Y(inst_ID2EX_reg_N73) );
  INVX1 U3351 ( .A(n4256), .Y(n4265) );
  INVX1 U3352 ( .A(n3387), .Y(inst_ID2EX_reg_N101) );
  INVX1 U3353 ( .A(n3162), .Y(inst_ID2EX_reg_N102) );
  INVX2 U3354 ( .A(n4426), .Y(n3805) );
  INVX4 U3355 ( .A(n4419), .Y(n4414) );
  INVX4 U3356 ( .A(n4753), .Y(n5002) );
  INVX4 U3357 ( .A(n4759), .Y(n4794) );
  INVX4 U3358 ( .A(n4877), .Y(n5119) );
  INVX4 U3359 ( .A(n2844), .Y(n3534) );
  INVX1 U3360 ( .A(n4080), .Y(n4084) );
  INVX1 U3361 ( .A(n4085), .Y(n4094) );
  INVX1 U3362 ( .A(n4212), .Y(n4099) );
  INVX1 U3363 ( .A(n4125), .Y(n4066) );
  INVX1 U3364 ( .A(n4194), .Y(n4195) );
  INVX1 U3365 ( .A(n4130), .Y(n4068) );
  INVX1 U3366 ( .A(n4058), .Y(n4061) );
  INVX1 U3367 ( .A(n4239), .Y(n4242) );
  INVX1 U3368 ( .A(n4215), .Y(n4217) );
  INVX1 U3369 ( .A(n4225), .Y(n4155) );
  INVX1 U3370 ( .A(n4236), .Y(n4237) );
  INVX1 U3371 ( .A(n4168), .Y(n4158) );
  INVX1 U3372 ( .A(n4226), .Y(n4235) );
  INVX1 U3373 ( .A(n2907), .Y(n2909) );
  INVX1 U3374 ( .A(n2928), .Y(n2929) );
  INVX1 U3375 ( .A(n4279), .Y(n3917) );
  INVX1 U3376 ( .A(n4440), .Y(n4441) );
  INVX1 U3377 ( .A(n4045), .Y(n3739) );
  INVX1 U3378 ( .A(n4254), .Y(n2972) );
  INVX1 U3379 ( .A(n3636), .Y(n3637) );
  INVX1 U3380 ( .A(n3925), .Y(n3918) );
  INVX1 U3381 ( .A(n4151), .Y(n4172) );
  INVX1 U3382 ( .A(n3985), .Y(n4174) );
  INVX1 U3383 ( .A(n3993), .Y(n4166) );
  INVX1 U3384 ( .A(n4063), .Y(n4136) );
  INVX1 U3385 ( .A(n4023), .Y(n4105) );
  INVX1 U3386 ( .A(n4399), .Y(n3643) );
  INVX1 U3387 ( .A(n4286), .Y(n4290) );
  INVX1 U3388 ( .A(n3928), .Y(n3930) );
  INVX1 U3389 ( .A(n5192), .Y(n5193) );
  INVX1 U3390 ( .A(n5189), .Y(n5190) );
  INVX1 U3391 ( .A(n3696), .Y(n5184) );
  INVX1 U3392 ( .A(n3685), .Y(n5182) );
  INVX1 U3393 ( .A(n4059), .Y(n4001) );
  INVX1 U3394 ( .A(n3652), .Y(n5176) );
  INVX1 U3395 ( .A(n5171), .Y(n5172) );
  INVX1 U3396 ( .A(n3506), .Y(n5169) );
  INVX1 U3397 ( .A(n3442), .Y(n5165) );
  INVX1 U3398 ( .A(n5162), .Y(n5163) );
  INVX1 U3399 ( .A(n5149), .Y(n5150) );
  INVX1 U3400 ( .A(n5144), .Y(n5145) );
  INVX1 U3401 ( .A(n5135), .Y(n5136) );
  INVX1 U3402 ( .A(n3434), .Y(n5124) );
  INVX1 U3403 ( .A(n5126), .Y(n5127) );
  INVX1 U3404 ( .A(n5231), .Y(n5232) );
  INVX1 U3405 ( .A(n4687), .Y(n4688) );
  INVX1 U3406 ( .A(n5518), .Y(n5516) );
  INVX1 U3407 ( .A(n3849), .Y(n4299) );
  INVX1 U3408 ( .A(n3850), .Y(n4293) );
  INVX1 U3409 ( .A(n2795), .Y(n3843) );
  INVX1 U3410 ( .A(n3960), .Y(n3965) );
  INVX1 U3411 ( .A(n3968), .Y(n3972) );
  INVX1 U3412 ( .A(n3975), .Y(n3979) );
  INVX1 U3413 ( .A(n3982), .Y(n3987) );
  INVX1 U3414 ( .A(n3990), .Y(n3995) );
  INVX1 U3415 ( .A(n3998), .Y(n4003) );
  INVX1 U3416 ( .A(n4006), .Y(n4010) );
  INVX1 U3417 ( .A(n4013), .Y(n4017) );
  INVX1 U3418 ( .A(n4020), .Y(n4025) );
  INVX1 U3419 ( .A(n4028), .Y(n4032) );
  INVX1 U3420 ( .A(n2795), .Y(n4312) );
  INVX1 U3421 ( .A(n2795), .Y(n3844) );
  INVX1 U3422 ( .A(n4327), .Y(n4328) );
  INVX1 U3423 ( .A(n3550), .Y(inst_ID2EX_reg_N68) );
  INVX1 U3424 ( .A(n3425), .Y(inst_ID2EX_reg_N67) );
  INVX1 U3425 ( .A(n3344), .Y(inst_ID2EX_reg_N99) );
  INVX1 U3426 ( .A(n3372), .Y(inst_ID2EX_reg_N98) );
  INVX1 U3427 ( .A(n3322), .Y(inst_ID2EX_reg_N65) );
  INVX1 U3428 ( .A(n3308), .Y(inst_ID2EX_reg_N97) );
  INVX1 U3429 ( .A(n3315), .Y(inst_ID2EX_reg_N96) );
  INVX1 U3430 ( .A(n3266), .Y(inst_ID2EX_reg_N63) );
  INVX1 U3431 ( .A(n3252), .Y(inst_ID2EX_reg_N95) );
  INVX1 U3432 ( .A(n3280), .Y(inst_ID2EX_reg_N94) );
  INVX1 U3433 ( .A(n3259), .Y(inst_ID2EX_reg_N61) );
  INVX1 U3434 ( .A(n3330), .Y(inst_ID2EX_reg_N60) );
  INVX1 U3435 ( .A(n3230), .Y(inst_ID2EX_reg_N92) );
  INVX1 U3436 ( .A(n3273), .Y(inst_ID2EX_reg_N59) );
  INVX1 U3437 ( .A(n3301), .Y(inst_ID2EX_reg_N58) );
  INVX1 U3438 ( .A(n3462), .Y(inst_ID2EX_reg_N90) );
  INVX1 U3439 ( .A(n3379), .Y(inst_ID2EX_reg_N57) );
  INVX1 U3440 ( .A(n3358), .Y(inst_ID2EX_reg_N56) );
  INVX1 U3441 ( .A(n3497), .Y(inst_ID2EX_reg_N88) );
  INVX1 U3442 ( .A(n2978), .Y(inst_EX2MEM_reg_N55) );
  INVX1 U3443 ( .A(n2992), .Y(inst_EX2MEM_reg_N54) );
  INVX1 U3444 ( .A(n3395), .Y(inst_ID2EX_reg_N86) );
  INVX1 U3445 ( .A(n3287), .Y(inst_ID2EX_reg_N53) );
  INVX1 U3446 ( .A(n3006), .Y(inst_EX2MEM_reg_N52) );
  INVX1 U3447 ( .A(n3558), .Y(inst_ID2EX_reg_N84) );
  INVX1 U3448 ( .A(n3476), .Y(inst_ID2EX_reg_N83) );
  INVX1 U3449 ( .A(n3094), .Y(inst_ID2EX_reg_N50) );
  INVX1 U3450 ( .A(n3409), .Y(inst_ID2EX_reg_N82) );
  INVX1 U3451 ( .A(n3469), .Y(inst_ID2EX_reg_N81) );
  INVX1 U3452 ( .A(n3013), .Y(inst_EX2MEM_reg_N48) );
  INVX1 U3453 ( .A(n3526), .Y(inst_ID2EX_reg_N80) );
  INVX1 U3454 ( .A(n3417), .Y(inst_ID2EX_reg_N79) );
  INVX1 U3455 ( .A(n3584), .Y(inst_EX2MEM_reg_N46) );
  INVX1 U3456 ( .A(n3577), .Y(inst_EX2MEM_reg_N45) );
  INVX1 U3457 ( .A(n3483), .Y(inst_ID2EX_reg_N77) );
  INVX1 U3458 ( .A(n3108), .Y(inst_ID2EX_reg_N44) );
  INVX1 U3459 ( .A(n3197), .Y(inst_EX2MEM_reg_N43) );
  INVX1 U3460 ( .A(n3533), .Y(inst_ID2EX_reg_N75) );
  INVX1 U3461 ( .A(n3204), .Y(inst_EX2MEM_reg_N42) );
  INVX1 U3462 ( .A(n3087), .Y(inst_ID2EX_reg_N39) );
  INVX1 U3463 ( .A(n3440), .Y(inst_ID2EX_reg_N71) );
  INVX1 U3464 ( .A(n3115), .Y(inst_ID2EX_reg_N40) );
  INVX1 U3465 ( .A(n3079), .Y(inst_ID2EX_reg_N41) );
  INVX1 U3466 ( .A(n3570), .Y(inst_ID2EX_reg_N69) );
  INVX1 U3467 ( .A(n3169), .Y(inst_ID2EX_reg_N70) );
  INVX1 U3468 ( .A(op_type_EX[1]), .Y(n2973) );
  BUFX2 U3469 ( .A(rst_n), .Y(n3066) );
  INVX2 U3470 ( .A(n3066), .Y(n5392) );
  INVX1 U3471 ( .A(alu_result_MEM[31]), .Y(n3769) );
  INVX1 U3472 ( .A(alu_result_MEM[27]), .Y(n3773) );
  INVX1 U3473 ( .A(alu_result_MEM[29]), .Y(n3771) );
  NAND3X1 U3474 ( .A(n3769), .B(n3773), .C(n3771), .Y(n2816) );
  NOR2X1 U3475 ( .A(alu_result_MEM[26]), .B(n2816), .Y(n2817) );
  INVX1 U3476 ( .A(alu_result_MEM[28]), .Y(n3772) );
  INVX1 U3477 ( .A(alu_result_MEM[30]), .Y(n3770) );
  NAND3X1 U3478 ( .A(n2817), .B(n3772), .C(n3770), .Y(n2834) );
  INVX1 U3479 ( .A(alu_result_MEM[23]), .Y(n3778) );
  INVX1 U3480 ( .A(alu_result_MEM[22]), .Y(n3779) );
  INVX1 U3481 ( .A(alu_result_MEM[18]), .Y(n3783) );
  NAND3X1 U3482 ( .A(n3778), .B(n3779), .C(n3783), .Y(n2818) );
  NOR2X1 U3483 ( .A(alu_result_MEM[19]), .B(n2818), .Y(n2819) );
  INVX1 U3484 ( .A(alu_result_MEM[20]), .Y(n3781) );
  INVX1 U3485 ( .A(alu_result_MEM[21]), .Y(n3780) );
  NAND3X1 U3486 ( .A(n2819), .B(n3781), .C(n3780), .Y(n2831) );
  INVX1 U3487 ( .A(alu_result_MEM[17]), .Y(n3784) );
  INVX1 U3488 ( .A(alu_result_MEM[10]), .Y(n3791) );
  INVX1 U3489 ( .A(alu_result_MEM[6]), .Y(n3795) );
  NAND3X1 U3490 ( .A(n3784), .B(n3791), .C(n3795), .Y(n2820) );
  NOR2X1 U3491 ( .A(alu_result_MEM[5]), .B(n2820), .Y(n2821) );
  INVX1 U3492 ( .A(alu_result_MEM[14]), .Y(n3787) );
  NAND3X1 U3493 ( .A(op_type_MEM[3]), .B(n2821), .C(n3787), .Y(n2828) );
  INVX1 U3494 ( .A(alu_result_MEM[0]), .Y(n4443) );
  INVX1 U3495 ( .A(alu_result_MEM[1]), .Y(n4434) );
  INVX1 U3496 ( .A(alu_result_MEM[2]), .Y(n4432) );
  NAND2X1 U3497 ( .A(n4434), .B(n4432), .Y(n4440) );
  NOR2X1 U3498 ( .A(n4443), .B(n4440), .Y(n4795) );
  INVX1 U3499 ( .A(alu_result_MEM[11]), .Y(n3790) );
  INVX1 U3500 ( .A(alu_result_MEM[12]), .Y(n3789) );
  NAND3X1 U3501 ( .A(n4795), .B(n3790), .C(n3789), .Y(n2825) );
  INVX1 U3502 ( .A(op_type_MEM[0]), .Y(n4430) );
  INVX1 U3503 ( .A(alu_result_MEM[3]), .Y(n3798) );
  INVX1 U3504 ( .A(op_type_MEM[1]), .Y(n3768) );
  INVX1 U3505 ( .A(op_type_MEM[2]), .Y(n4429) );
  NAND2X1 U3506 ( .A(n3768), .B(n4429), .Y(n2845) );
  INVX1 U3507 ( .A(alu_result_MEM[8]), .Y(n3793) );
  INVX1 U3508 ( .A(alu_result_MEM[25]), .Y(n3776) );
  INVX1 U3509 ( .A(alu_result_MEM[24]), .Y(n3777) );
  NAND3X1 U3510 ( .A(n3793), .B(n3776), .C(n3777), .Y(n2822) );
  NOR2X1 U3511 ( .A(n2845), .B(n2822), .Y(n2823) );
  NAND3X1 U3512 ( .A(n4430), .B(n3798), .C(n2823), .Y(n2824) );
  NOR2X1 U3513 ( .A(n2825), .B(n2824), .Y(n2826) );
  INVX1 U3514 ( .A(alu_result_MEM[4]), .Y(n3797) );
  INVX1 U3515 ( .A(alu_result_MEM[15]), .Y(n3786) );
  NAND3X1 U3516 ( .A(n2826), .B(n3797), .C(n3786), .Y(n2827) );
  NOR2X1 U3517 ( .A(n2828), .B(n2827), .Y(n2829) );
  INVX1 U3518 ( .A(alu_result_MEM[16]), .Y(n3785) );
  INVX1 U3519 ( .A(alu_result_MEM[13]), .Y(n3788) );
  NAND3X1 U3520 ( .A(n2829), .B(n3785), .C(n3788), .Y(n2830) );
  NOR2X1 U3521 ( .A(n2831), .B(n2830), .Y(n2832) );
  INVX1 U3522 ( .A(alu_result_MEM[7]), .Y(n3794) );
  INVX1 U3523 ( .A(alu_result_MEM[9]), .Y(n3792) );
  NAND3X1 U3524 ( .A(n2832), .B(n3794), .C(n3792), .Y(n2833) );
  NOR2X1 U3525 ( .A(n2834), .B(n2833), .Y(n3634) );
  NAND2X1 U3526 ( .A(op_type_MEM[3]), .B(op_type_MEM[0]), .Y(n2835) );
  NOR2X1 U3527 ( .A(n2845), .B(n2835), .Y(n3636) );
  NOR2X1 U3528 ( .A(n3634), .B(n3636), .Y(n4616) );
  AND2X2 U3529 ( .A(n2815), .B(n4616), .Y(n4426) );
  NOR2X1 U3530 ( .A(n2973), .B(n3774), .Y(inst_EX2MEM_reg_N4) );
  INVX1 U3531 ( .A(op_type_EX[2]), .Y(n4193) );
  NOR2X1 U3532 ( .A(n4193), .B(n2809), .Y(inst_EX2MEM_reg_N5) );
  INVX1 U3533 ( .A(op_type_EX[3]), .Y(n3804) );
  NAND2X1 U3534 ( .A(op_type_EX[2]), .B(n3804), .Y(n4183) );
  INVX1 U3535 ( .A(n4183), .Y(n2836) );
  NAND2X1 U3536 ( .A(n2836), .B(op_type_EX[1]), .Y(n3045) );
  NOR2X1 U3537 ( .A(op_type_EX[2]), .B(op_type_EX[3]), .Y(n2837) );
  NAND3X1 U3538 ( .A(op_type_EX[0]), .B(n2973), .C(n2837), .Y(n2840) );
  NOR2X1 U3539 ( .A(op_type_EX[3]), .B(op_type_EX[0]), .Y(n2971) );
  NAND2X1 U3540 ( .A(n2971), .B(op_type_EX[1]), .Y(n2838) );
  INVX4 U3541 ( .A(n2839), .Y(n4259) );
  NAND3X1 U3542 ( .A(n3045), .B(n2840), .C(n2839), .Y(n2841) );
  NAND2X1 U3543 ( .A(n2841), .B(n4426), .Y(n4033) );
  INVX1 U3544 ( .A(op_type_WB[2]), .Y(n2842) );
  NOR2X1 U3545 ( .A(op_type_WB[0]), .B(n2842), .Y(n2858) );
  NAND2X1 U3546 ( .A(n2858), .B(op_type_WB[1]), .Y(n2843) );
  MUX2X1 U3547 ( .B(alu_result_WB[16]), .A(mem_read_data_WB[16]), .S(n3534), 
        .Y(n3506) );
  NAND3X1 U3548 ( .A(op_type_MEM[1]), .B(op_type_MEM[0]), .C(op_type_MEM[2]), 
        .Y(n3592) );
  OAI21X1 U3549 ( .A(op_type_MEM[0]), .B(n2845), .C(n3592), .Y(n2846) );
  NOR2X1 U3550 ( .A(op_type_MEM[3]), .B(n2846), .Y(n2875) );
  INVX1 U3551 ( .A(reg_write_address_MEM[3]), .Y(n3800) );
  INVX1 U3552 ( .A(read_register_1_EX[0]), .Y(n3749) );
  INVX1 U3553 ( .A(reg_write_address_MEM[0]), .Y(n3803) );
  AOI22X1 U3554 ( .A(reg_write_address_MEM[0]), .B(n3749), .C(
        read_register_1_EX[0]), .D(n3803), .Y(n2847) );
  OAI21X1 U3555 ( .A(read_register_1_EX[3]), .B(n3800), .C(n2847), .Y(n2848)
         );
  AOI21X1 U3556 ( .A(read_register_1_EX[3]), .B(n3800), .C(n2848), .Y(n2854)
         );
  INVX1 U3557 ( .A(reg_write_address_MEM[2]), .Y(n3801) );
  INVX1 U3558 ( .A(read_register_1_EX[4]), .Y(n3745) );
  INVX1 U3559 ( .A(read_register_1_EX[1]), .Y(n3748) );
  INVX1 U3560 ( .A(reg_write_address_MEM[1]), .Y(n3802) );
  AOI22X1 U3561 ( .A(reg_write_address_MEM[1]), .B(n3748), .C(
        read_register_1_EX[1]), .D(n3802), .Y(n2849) );
  OAI21X1 U3562 ( .A(reg_write_address_MEM[4]), .B(n3745), .C(n2849), .Y(n2850) );
  AOI21X1 U3563 ( .A(reg_write_address_MEM[4]), .B(n3745), .C(n2850), .Y(n2851) );
  OAI21X1 U3564 ( .A(read_register_1_EX[2]), .B(n3801), .C(n2851), .Y(n2852)
         );
  AOI21X1 U3565 ( .A(read_register_1_EX[2]), .B(n3801), .C(n2852), .Y(n2853)
         );
  NAND3X1 U3566 ( .A(n2875), .B(n2854), .C(n2853), .Y(n2868) );
  INVX1 U3567 ( .A(reg_write_address_WB[4]), .Y(n3137) );
  INVX1 U3568 ( .A(read_register_1_EX[2]), .Y(n3747) );
  INVX1 U3569 ( .A(reg_write_address_WB[0]), .Y(n5201) );
  AOI22X1 U3570 ( .A(reg_write_address_WB[0]), .B(n3749), .C(
        read_register_1_EX[0]), .D(n5201), .Y(n2855) );
  OAI21X1 U3571 ( .A(reg_write_address_WB[2]), .B(n3747), .C(n2855), .Y(n2865)
         );
  INVX1 U3572 ( .A(reg_write_address_WB[2]), .Y(n5391) );
  INVX1 U3573 ( .A(reg_write_address_WB[3]), .Y(n3139) );
  INVX1 U3574 ( .A(reg_write_address_WB[1]), .Y(n5428) );
  AOI22X1 U3575 ( .A(reg_write_address_WB[1]), .B(n3748), .C(
        read_register_1_EX[1]), .D(n5428), .Y(n2856) );
  OAI21X1 U3576 ( .A(read_register_1_EX[3]), .B(n3139), .C(n2856), .Y(n2862)
         );
  INVX1 U3577 ( .A(read_register_1_EX[3]), .Y(n3746) );
  NAND2X1 U3578 ( .A(op_type_WB[2]), .B(op_type_WB[1]), .Y(n2857) );
  OAI21X1 U3579 ( .A(op_type_WB[1]), .B(op_type_WB[0]), .C(n2857), .Y(n2860)
         );
  INVX1 U3580 ( .A(n2858), .Y(n2859) );
  AOI21X1 U3581 ( .A(n2860), .B(n2859), .C(op_type_WB[3]), .Y(n5202) );
  OAI21X1 U3582 ( .A(reg_write_address_WB[3]), .B(n3746), .C(n5202), .Y(n2861)
         );
  NOR2X1 U3583 ( .A(n2862), .B(n2861), .Y(n2863) );
  OAI21X1 U3584 ( .A(read_register_1_EX[2]), .B(n5391), .C(n2863), .Y(n2864)
         );
  NOR2X1 U3585 ( .A(n2865), .B(n2864), .Y(n2866) );
  OAI21X1 U3586 ( .A(read_register_1_EX[4]), .B(n3137), .C(n2866), .Y(n2867)
         );
  AOI21X1 U3587 ( .A(read_register_1_EX[4]), .B(n3137), .C(n2867), .Y(n2869)
         );
  NAND2X1 U3588 ( .A(n2868), .B(n2869), .Y(n3733) );
  INVX4 U3589 ( .A(n2870), .Y(n3947) );
  AOI22X1 U3590 ( .A(reg_read_data_1_EX[16]), .B(n3947), .C(alu_result_MEM[16]), .D(n2814), .Y(n2871) );
  OAI21X1 U3591 ( .A(n3506), .B(n3733), .C(n2871), .Y(n4112) );
  BUFX2 U3592 ( .A(n3045), .Y(n2965) );
  INVX1 U3593 ( .A(n2965), .Y(n2872) );
  INVX1 U3594 ( .A(jump_inst_addr_EX[15]), .Y(n4419) );
  NAND2X1 U3595 ( .A(n2872), .B(n4414), .Y(n3943) );
  INVX1 U3596 ( .A(read_register_2_EX[4]), .Y(n3750) );
  INVX1 U3597 ( .A(read_register_2_EX[1]), .Y(n3753) );
  AOI22X1 U3598 ( .A(read_register_2_EX[1]), .B(n3802), .C(
        reg_write_address_MEM[1]), .D(n3753), .Y(n2873) );
  OAI21X1 U3599 ( .A(read_register_2_EX[3]), .B(n3800), .C(n2873), .Y(n2880)
         );
  INVX1 U3600 ( .A(read_register_2_EX[3]), .Y(n3751) );
  INVX1 U3601 ( .A(read_register_2_EX[2]), .Y(n3752) );
  INVX1 U3602 ( .A(read_register_2_EX[0]), .Y(n3754) );
  AOI22X1 U3603 ( .A(read_register_2_EX[0]), .B(n3803), .C(
        reg_write_address_MEM[0]), .D(n3754), .Y(n2874) );
  OAI21X1 U3604 ( .A(reg_write_address_MEM[2]), .B(n3752), .C(n2874), .Y(n2877) );
  OAI21X1 U3605 ( .A(read_register_2_EX[2]), .B(n3801), .C(n2875), .Y(n2876)
         );
  NOR2X1 U3606 ( .A(n2877), .B(n2876), .Y(n2878) );
  OAI21X1 U3607 ( .A(reg_write_address_MEM[3]), .B(n3751), .C(n2878), .Y(n2879) );
  NOR2X1 U3608 ( .A(n2880), .B(n2879), .Y(n2881) );
  OAI21X1 U3609 ( .A(reg_write_address_MEM[4]), .B(n3750), .C(n2881), .Y(n2882) );
  AOI21X1 U3610 ( .A(reg_write_address_MEM[4]), .B(n3750), .C(n2882), .Y(n2892) );
  NAND2X1 U3611 ( .A(n2892), .B(n2965), .Y(n3720) );
  INVX4 U3612 ( .A(n3720), .Y(n3942) );
  AOI22X1 U3613 ( .A(read_register_2_EX[4]), .B(n3137), .C(
        reg_write_address_WB[4]), .D(n3750), .Y(n2883) );
  OAI21X1 U3614 ( .A(read_register_2_EX[2]), .B(n5391), .C(n2883), .Y(n2889)
         );
  AOI22X1 U3615 ( .A(read_register_2_EX[0]), .B(n5201), .C(
        reg_write_address_WB[0]), .D(n3754), .Y(n2884) );
  OAI21X1 U3616 ( .A(reg_write_address_WB[1]), .B(n3753), .C(n2884), .Y(n2886)
         );
  OAI21X1 U3617 ( .A(read_register_2_EX[1]), .B(n5428), .C(n5202), .Y(n2885)
         );
  NOR2X1 U3618 ( .A(n2886), .B(n2885), .Y(n2887) );
  OAI21X1 U3619 ( .A(reg_write_address_WB[2]), .B(n3752), .C(n2887), .Y(n2888)
         );
  NOR2X1 U3620 ( .A(n2889), .B(n2888), .Y(n2890) );
  OAI21X1 U3621 ( .A(read_register_2_EX[3]), .B(n3139), .C(n2890), .Y(n2891)
         );
  AOI21X1 U3622 ( .A(read_register_2_EX[3]), .B(n3139), .C(n2891), .Y(n2896)
         );
  INVX1 U3623 ( .A(n2892), .Y(n2893) );
  NAND2X1 U3624 ( .A(n2965), .B(n2893), .Y(n2897) );
  INVX4 U3625 ( .A(n2894), .Y(n3941) );
  AOI22X1 U3626 ( .A(alu_result_MEM[16]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[16]), .Y(n2895) );
  AND2X2 U3627 ( .A(n3943), .B(n2895), .Y(n2900) );
  INVX1 U3628 ( .A(n2896), .Y(n2898) );
  NOR2X1 U3629 ( .A(n2898), .B(n2897), .Y(n3946) );
  NAND2X1 U3630 ( .A(n5169), .B(n3946), .Y(n2899) );
  NAND2X1 U3631 ( .A(n2900), .B(n2899), .Y(n4130) );
  XOR2X1 U3632 ( .A(n4259), .B(n4130), .Y(n3663) );
  MUX2X1 U3633 ( .B(alu_result_WB[15]), .A(mem_read_data_WB[15]), .S(n3534), 
        .Y(n3389) );
  AOI22X1 U3634 ( .A(reg_read_data_1_EX[15]), .B(n3947), .C(alu_result_MEM[15]), .D(n2814), .Y(n2902) );
  OAI21X1 U3635 ( .A(n3389), .B(n2901), .C(n2902), .Y(n4124) );
  AOI22X1 U3636 ( .A(alu_result_MEM[15]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[15]), .Y(n2904) );
  NAND2X1 U3637 ( .A(n5167), .B(n3946), .Y(n2903) );
  NAND3X1 U3638 ( .A(n3943), .B(n2904), .C(n2903), .Y(n4125) );
  XOR2X1 U3639 ( .A(n4259), .B(n4125), .Y(n2987) );
  MUX2X1 U3640 ( .B(alu_result_WB[14]), .A(mem_read_data_WB[14]), .S(n3534), 
        .Y(n3442) );
  AOI22X1 U3641 ( .A(reg_read_data_1_EX[14]), .B(n3947), .C(alu_result_MEM[14]), .D(n2814), .Y(n2905) );
  OAI21X1 U3642 ( .A(n3442), .B(n2901), .C(n2905), .Y(n4120) );
  INVX1 U3643 ( .A(jump_inst_addr_EX[14]), .Y(n3755) );
  AOI22X1 U3644 ( .A(alu_result_MEM[14]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[14]), .Y(n2906) );
  OAI21X1 U3645 ( .A(n2965), .B(n3755), .C(n2906), .Y(n2907) );
  NAND2X1 U3646 ( .A(n5165), .B(n3946), .Y(n2908) );
  NAND2X1 U3647 ( .A(n2909), .B(n2908), .Y(n4065) );
  XOR2X1 U3648 ( .A(n4259), .B(n4065), .Y(n2980) );
  MUX2X1 U3649 ( .B(alu_result_WB[13]), .A(mem_read_data_WB[13]), .S(n3534), 
        .Y(n5162) );
  AOI22X1 U3650 ( .A(reg_read_data_1_EX[13]), .B(n3947), .C(alu_result_MEM[13]), .D(n2814), .Y(n2910) );
  OAI21X1 U3651 ( .A(n5162), .B(n2901), .C(n2910), .Y(n4114) );
  INVX1 U3652 ( .A(jump_inst_addr_EX[13]), .Y(n3756) );
  AOI22X1 U3653 ( .A(alu_result_MEM[13]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[13]), .Y(n2911) );
  OAI21X1 U3654 ( .A(n3045), .B(n3756), .C(n2911), .Y(n2912) );
  OAI21X1 U3655 ( .A(n5162), .B(n3736), .C(n2913), .Y(n4117) );
  XOR2X1 U3656 ( .A(n4259), .B(n4117), .Y(n3001) );
  MUX2X1 U3657 ( .B(alu_result_WB[12]), .A(mem_read_data_WB[12]), .S(n3534), 
        .Y(n5159) );
  AOI22X1 U3658 ( .A(reg_read_data_1_EX[12]), .B(n3947), .C(alu_result_MEM[12]), .D(n2814), .Y(n2914) );
  OAI21X1 U3659 ( .A(n5159), .B(n2901), .C(n2914), .Y(n4110) );
  INVX1 U3660 ( .A(jump_inst_addr_EX[12]), .Y(n4375) );
  AOI22X1 U3661 ( .A(alu_result_MEM[12]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[12]), .Y(n2915) );
  OAI21X1 U3662 ( .A(n2965), .B(n4375), .C(n2915), .Y(n2916) );
  OAI21X1 U3663 ( .A(n5159), .B(n3736), .C(n2917), .Y(n4115) );
  XOR2X1 U3664 ( .A(n4259), .B(n4115), .Y(n2994) );
  MUX2X1 U3665 ( .B(alu_result_WB[11]), .A(mem_read_data_WB[11]), .S(n3534), 
        .Y(n5156) );
  AOI22X1 U3666 ( .A(reg_read_data_1_EX[11]), .B(n3947), .C(alu_result_MEM[11]), .D(n2814), .Y(n2918) );
  OAI21X1 U3667 ( .A(n5156), .B(n2901), .C(n2918), .Y(n4023) );
  INVX1 U3668 ( .A(jump_inst_addr_EX[11]), .Y(n3757) );
  AOI22X1 U3669 ( .A(alu_result_MEM[11]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[11]), .Y(n2919) );
  OAI21X1 U3670 ( .A(n3045), .B(n3757), .C(n2919), .Y(n2920) );
  OAI21X1 U3671 ( .A(n5156), .B(n3736), .C(n2921), .Y(n4104) );
  XOR2X1 U3672 ( .A(n4259), .B(n4104), .Y(n4019) );
  MUX2X1 U3673 ( .B(alu_result_WB[10]), .A(mem_read_data_WB[10]), .S(n3534), 
        .Y(n5152) );
  AOI22X1 U3674 ( .A(reg_read_data_1_EX[10]), .B(n3947), .C(alu_result_MEM[10]), .D(n2814), .Y(n2922) );
  OAI21X1 U3675 ( .A(n5152), .B(n2901), .C(n2922), .Y(n4101) );
  INVX1 U3676 ( .A(jump_inst_addr_EX[10]), .Y(n3758) );
  AOI22X1 U3677 ( .A(alu_result_MEM[10]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[10]), .Y(n2923) );
  OAI21X1 U3678 ( .A(n2965), .B(n3758), .C(n2923), .Y(n2924) );
  OAI21X1 U3679 ( .A(n5152), .B(n3736), .C(n2925), .Y(n4106) );
  XOR2X1 U3680 ( .A(n4259), .B(n4106), .Y(n3015) );
  MUX2X1 U3681 ( .B(alu_result_WB[9]), .A(mem_read_data_WB[9]), .S(n3534), .Y(
        n5149) );
  AOI22X1 U3682 ( .A(reg_read_data_1_EX[9]), .B(n3947), .C(alu_result_MEM[9]), 
        .D(n2814), .Y(n2926) );
  OAI21X1 U3683 ( .A(n5149), .B(n2901), .C(n2926), .Y(n4096) );
  INVX1 U3684 ( .A(jump_inst_addr_EX[9]), .Y(n4367) );
  AOI22X1 U3685 ( .A(alu_result_MEM[9]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[9]), .Y(n2927) );
  OAI21X1 U3686 ( .A(n3045), .B(n4367), .C(n2927), .Y(n2928) );
  OAI21X1 U3687 ( .A(n5149), .B(n3736), .C(n2929), .Y(n4102) );
  XOR2X1 U3688 ( .A(n4259), .B(n4102), .Y(n3008) );
  MUX2X1 U3689 ( .B(alu_result_WB[8]), .A(mem_read_data_WB[8]), .S(n3534), .Y(
        n3411) );
  AOI22X1 U3690 ( .A(reg_read_data_1_EX[8]), .B(n3947), .C(alu_result_MEM[8]), 
        .D(n2814), .Y(n2930) );
  OAI21X1 U3691 ( .A(n3411), .B(n2901), .C(n2930), .Y(n4095) );
  INVX1 U3692 ( .A(jump_inst_addr_EX[8]), .Y(n3759) );
  AOI22X1 U3693 ( .A(alu_result_MEM[8]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[8]), .Y(n2931) );
  OAI21X1 U3694 ( .A(n2965), .B(n3759), .C(n2931), .Y(n2932) );
  NAND2X1 U3695 ( .A(n5147), .B(n3946), .Y(n2933) );
  NAND2X1 U3696 ( .A(n2934), .B(n2933), .Y(n4098) );
  XOR2X1 U3697 ( .A(n4259), .B(n4098), .Y(n3586) );
  MUX2X1 U3698 ( .B(alu_result_WB[7]), .A(mem_read_data_WB[7]), .S(n3534), .Y(
        n5144) );
  AOI22X1 U3699 ( .A(reg_read_data_1_EX[7]), .B(n3947), .C(alu_result_MEM[7]), 
        .D(n2814), .Y(n2935) );
  OAI21X1 U3700 ( .A(n5144), .B(n2901), .C(n2935), .Y(n4089) );
  INVX1 U3701 ( .A(jump_inst_addr_EX[7]), .Y(n3760) );
  AOI22X1 U3702 ( .A(alu_result_MEM[7]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[7]), .Y(n2936) );
  OAI21X1 U3703 ( .A(n3045), .B(n3760), .C(n2936), .Y(n2937) );
  OAI21X1 U3704 ( .A(n5144), .B(n3736), .C(n2938), .Y(n4090) );
  XOR2X1 U3705 ( .A(n4259), .B(n4090), .Y(n3579) );
  MUX2X1 U3706 ( .B(alu_result_WB[6]), .A(mem_read_data_WB[6]), .S(n3534), .Y(
        n5141) );
  AOI22X1 U3707 ( .A(reg_read_data_1_EX[6]), .B(n3947), .C(alu_result_MEM[6]), 
        .D(n2814), .Y(n2939) );
  OAI21X1 U3708 ( .A(n5141), .B(n2901), .C(n2939), .Y(n4086) );
  INVX1 U3709 ( .A(jump_inst_addr_EX[6]), .Y(n3761) );
  AOI22X1 U3710 ( .A(alu_result_MEM[6]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[6]), .Y(n2940) );
  OAI21X1 U3711 ( .A(n2965), .B(n3761), .C(n2940), .Y(n2941) );
  OAI21X1 U3712 ( .A(n5141), .B(n3736), .C(n2942), .Y(n4092) );
  XOR2X1 U3713 ( .A(n4259), .B(n4092), .Y(n3572) );
  MUX2X1 U3714 ( .B(alu_result_WB[5]), .A(mem_read_data_WB[5]), .S(n3534), .Y(
        n5138) );
  AOI22X1 U3715 ( .A(reg_read_data_1_EX[5]), .B(n3947), .C(alu_result_MEM[5]), 
        .D(n2814), .Y(n2943) );
  OAI21X1 U3716 ( .A(n5138), .B(n2901), .C(n2943), .Y(n4081) );
  INVX1 U3717 ( .A(jump_inst_addr_EX[5]), .Y(n3762) );
  AOI22X1 U3718 ( .A(n3941), .B(reg_read_data_2_EX[5]), .C(alu_result_MEM[5]), 
        .D(n3942), .Y(n2944) );
  OAI21X1 U3719 ( .A(n3045), .B(n3762), .C(n2944), .Y(n2945) );
  INVX1 U3720 ( .A(n2945), .Y(n2946) );
  OAI21X1 U3721 ( .A(n5138), .B(n3736), .C(n2946), .Y(n4087) );
  XOR2X1 U3722 ( .A(n4259), .B(n4087), .Y(n4027) );
  MUX2X1 U3723 ( .B(alu_result_WB[4]), .A(mem_read_data_WB[4]), .S(n3534), .Y(
        n5135) );
  AOI22X1 U3724 ( .A(reg_read_data_1_EX[4]), .B(n3947), .C(alu_result_MEM[4]), 
        .D(n2814), .Y(n2947) );
  OAI21X1 U3725 ( .A(n5135), .B(n2901), .C(n2947), .Y(n4071) );
  INVX1 U3726 ( .A(jump_inst_addr_EX[4]), .Y(n3763) );
  AOI22X1 U3727 ( .A(alu_result_MEM[4]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[4]), .Y(n2948) );
  OAI21X1 U3728 ( .A(n2965), .B(n3763), .C(n2948), .Y(n2949) );
  INVX1 U3729 ( .A(n2949), .Y(n2950) );
  OAI21X1 U3730 ( .A(n5135), .B(n3736), .C(n2950), .Y(n4083) );
  XOR2X1 U3731 ( .A(n4259), .B(n4083), .Y(n3192) );
  MUX2X1 U3732 ( .B(alu_result_WB[3]), .A(mem_read_data_WB[3]), .S(n3534), .Y(
        n5132) );
  AOI22X1 U3733 ( .A(reg_read_data_1_EX[3]), .B(n3947), .C(alu_result_MEM[3]), 
        .D(n2814), .Y(n2951) );
  OAI21X1 U3734 ( .A(n5132), .B(n2901), .C(n2951), .Y(n4072) );
  INVX1 U3735 ( .A(jump_inst_addr_EX[3]), .Y(n3764) );
  AOI22X1 U3736 ( .A(alu_result_MEM[3]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[3]), .Y(n2952) );
  OAI21X1 U3737 ( .A(n2965), .B(n3764), .C(n2952), .Y(n2953) );
  INVX1 U3738 ( .A(n2953), .Y(n2954) );
  OAI21X1 U3739 ( .A(n5132), .B(n3736), .C(n2954), .Y(n4077) );
  XOR2X1 U3740 ( .A(n4259), .B(n4077), .Y(n3199) );
  MUX2X1 U3741 ( .B(alu_result_WB[2]), .A(mem_read_data_WB[2]), .S(n3534), .Y(
        n5129) );
  AOI22X1 U3742 ( .A(reg_read_data_1_EX[2]), .B(n3947), .C(alu_result_MEM[2]), 
        .D(n2814), .Y(n2955) );
  OAI21X1 U3743 ( .A(n5129), .B(n2901), .C(n2955), .Y(n4039) );
  INVX1 U3744 ( .A(jump_inst_addr_EX[2]), .Y(n3765) );
  AOI22X1 U3745 ( .A(n3941), .B(reg_read_data_2_EX[2]), .C(alu_result_MEM[2]), 
        .D(n3942), .Y(n2956) );
  OAI21X1 U3746 ( .A(n2965), .B(n3765), .C(n2956), .Y(n2957) );
  INVX1 U3747 ( .A(n2957), .Y(n2958) );
  OAI21X1 U3748 ( .A(n5129), .B(n3736), .C(n2958), .Y(n4075) );
  XOR2X1 U3749 ( .A(n4259), .B(n4075), .Y(n4035) );
  MUX2X1 U3750 ( .B(alu_result_WB[1]), .A(mem_read_data_WB[1]), .S(n3534), .Y(
        n5126) );
  AOI22X1 U3751 ( .A(reg_read_data_1_EX[1]), .B(n3947), .C(alu_result_MEM[1]), 
        .D(n2814), .Y(n2959) );
  OAI21X1 U3752 ( .A(n5126), .B(n2901), .C(n2959), .Y(n4201) );
  INVX1 U3753 ( .A(jump_inst_addr_EX[1]), .Y(n3766) );
  AOI22X1 U3754 ( .A(n3941), .B(reg_read_data_2_EX[1]), .C(alu_result_MEM[1]), 
        .D(n3942), .Y(n2960) );
  OAI21X1 U3755 ( .A(n2965), .B(n3766), .C(n2960), .Y(n2961) );
  INVX1 U3756 ( .A(n2961), .Y(n2962) );
  OAI21X1 U3757 ( .A(n5126), .B(n3736), .C(n2962), .Y(n4191) );
  XOR2X1 U3758 ( .A(n4259), .B(n4191), .Y(n4043) );
  MUX2X1 U3759 ( .B(alu_result_WB[0]), .A(mem_read_data_WB[0]), .S(n3534), .Y(
        n3434) );
  AOI22X1 U3760 ( .A(reg_read_data_1_EX[0]), .B(n3947), .C(alu_result_MEM[0]), 
        .D(n2814), .Y(n2963) );
  OAI21X1 U3761 ( .A(n3434), .B(n2901), .C(n2963), .Y(n4258) );
  INVX1 U3762 ( .A(jump_inst_addr_EX[0]), .Y(n4332) );
  AOI22X1 U3763 ( .A(n3942), .B(alu_result_MEM[0]), .C(n3941), .D(
        reg_read_data_2_EX[0]), .Y(n2964) );
  OAI21X1 U3764 ( .A(n2965), .B(n4332), .C(n2964), .Y(n2966) );
  INVX1 U3765 ( .A(n2966), .Y(n2968) );
  NAND2X1 U3766 ( .A(n5124), .B(n3946), .Y(n2967) );
  NAND2X1 U3767 ( .A(n2968), .B(n2967), .Y(n4186) );
  XOR2X1 U3768 ( .A(n4259), .B(n4186), .Y(n4257) );
  NAND2X1 U3769 ( .A(n4112), .B(n4130), .Y(n2975) );
  NAND3X1 U3770 ( .A(op_type_EX[0]), .B(n4193), .C(n3804), .Y(n2969) );
  NAND2X1 U3771 ( .A(n2970), .B(inst_EX2MEM_reg_N4), .Y(n4047) );
  BUFX2 U3772 ( .A(n4047), .Y(n3953) );
  NAND2X1 U3773 ( .A(n2971), .B(inst_EX2MEM_reg_N5), .Y(n4254) );
  NAND2X1 U3774 ( .A(n2973), .B(n2972), .Y(n4045) );
  OAI21X1 U3775 ( .A(n4112), .B(n4130), .C(n3739), .Y(n2974) );
  OAI21X1 U3776 ( .A(n2975), .B(n3953), .C(n2974), .Y(n2976) );
  AOI21X1 U3777 ( .A(n4263), .B(n2977), .C(n2976), .Y(n2978) );
  FAX1 U3778 ( .A(n4120), .B(n2980), .C(n2979), .YC(n2986), .YS(n2984) );
  NAND2X1 U3779 ( .A(n4120), .B(n4065), .Y(n2982) );
  OAI21X1 U3780 ( .A(n4065), .B(n4120), .C(n3739), .Y(n2981) );
  OAI21X1 U3781 ( .A(n2982), .B(n3953), .C(n2981), .Y(n2983) );
  AOI21X1 U3782 ( .A(n4263), .B(n2984), .C(n2983), .Y(n2985) );
  FAX1 U3783 ( .A(n4124), .B(n2987), .C(n2986), .YC(n3662), .YS(n2991) );
  NAND2X1 U3784 ( .A(n4124), .B(n4125), .Y(n2989) );
  OAI21X1 U3785 ( .A(n4125), .B(n4124), .C(n3739), .Y(n2988) );
  OAI21X1 U3786 ( .A(n2989), .B(n4047), .C(n2988), .Y(n2990) );
  AOI21X1 U3787 ( .A(n4263), .B(n2991), .C(n2990), .Y(n2992) );
  FAX1 U3788 ( .A(n4110), .B(n2994), .C(n2993), .YC(n3000), .YS(n2998) );
  NAND2X1 U3789 ( .A(n4110), .B(n4115), .Y(n2996) );
  OAI21X1 U3790 ( .A(n4115), .B(n4110), .C(n3739), .Y(n2995) );
  OAI21X1 U3791 ( .A(n2996), .B(n4047), .C(n2995), .Y(n2997) );
  AOI21X1 U3792 ( .A(n4263), .B(n2998), .C(n2997), .Y(n2999) );
  FAX1 U3793 ( .A(n4114), .B(n3001), .C(n3000), .YC(n2979), .YS(n3005) );
  NAND2X1 U3794 ( .A(n4114), .B(n4117), .Y(n3003) );
  OAI21X1 U3795 ( .A(n4117), .B(n4114), .C(n3739), .Y(n3002) );
  OAI21X1 U3796 ( .A(n3003), .B(n4047), .C(n3002), .Y(n3004) );
  AOI21X1 U3797 ( .A(n4263), .B(n3005), .C(n3004), .Y(n3006) );
  FAX1 U3798 ( .A(n4096), .B(n3008), .C(n3007), .YC(n3014), .YS(n3012) );
  NAND2X1 U3799 ( .A(n4096), .B(n4102), .Y(n3010) );
  OAI21X1 U3800 ( .A(n4102), .B(n4096), .C(n3739), .Y(n3009) );
  OAI21X1 U3801 ( .A(n3010), .B(n4047), .C(n3009), .Y(n3011) );
  AOI21X1 U3802 ( .A(n4263), .B(n3012), .C(n3011), .Y(n3013) );
  FAX1 U3803 ( .A(n4101), .B(n3015), .C(n3014), .YC(n4018), .YS(n3019) );
  NAND2X1 U3804 ( .A(n4101), .B(n4106), .Y(n3017) );
  OAI21X1 U3805 ( .A(n4106), .B(n4101), .C(n3739), .Y(n3016) );
  OAI21X1 U3806 ( .A(n3017), .B(n3953), .C(n3016), .Y(n3018) );
  AOI21X1 U3807 ( .A(n4263), .B(n3019), .C(n3018), .Y(n3020) );
  INVX1 U3808 ( .A(instruction_ID[24]), .Y(n4634) );
  INVX1 U3809 ( .A(instruction_ID[22]), .Y(n4638) );
  AOI22X1 U3810 ( .A(reg_write_address_WB[1]), .B(instruction_ID[22]), .C(
        n4638), .D(n5428), .Y(n3026) );
  INVX1 U3811 ( .A(instruction_ID[25]), .Y(n4632) );
  AOI22X1 U3812 ( .A(reg_write_address_WB[4]), .B(n4632), .C(
        instruction_ID[25]), .D(n3137), .Y(n3021) );
  OAI21X1 U3813 ( .A(instruction_ID[23]), .B(n5391), .C(n3021), .Y(n3023) );
  INVX1 U3814 ( .A(instruction_ID[23]), .Y(n4636) );
  OAI21X1 U3815 ( .A(reg_write_address_WB[2]), .B(n4636), .C(n5202), .Y(n3022)
         );
  NOR2X1 U3816 ( .A(n3023), .B(n3022), .Y(n3024) );
  OAI21X1 U3817 ( .A(instruction_ID[24]), .B(n3139), .C(n3024), .Y(n3025) );
  NOR2X1 U3818 ( .A(n3026), .B(n3025), .Y(n3027) );
  OAI21X1 U3819 ( .A(reg_write_address_WB[3]), .B(n4634), .C(n3027), .Y(n3028)
         );
  AOI21X1 U3820 ( .A(n5201), .B(instruction_ID[21]), .C(n3028), .Y(n3029) );
  OAI21X1 U3821 ( .A(n5201), .B(instruction_ID[21]), .C(n3029), .Y(n3561) );
  INVX1 U3822 ( .A(instruction_ID[21]), .Y(n4640) );
  NAND2X1 U3823 ( .A(n4640), .B(n3030), .Y(n3040) );
  NAND2X1 U3824 ( .A(instruction_ID[23]), .B(n4638), .Y(n3036) );
  NOR2X1 U3825 ( .A(n3040), .B(n3036), .Y(n3564) );
  NAND2X1 U3826 ( .A(n4636), .B(n4638), .Y(n3039) );
  NAND2X1 U3827 ( .A(instruction_ID[21]), .B(n3030), .Y(n3035) );
  NOR2X1 U3828 ( .A(n3039), .B(n3035), .Y(n3563) );
  AOI22X1 U3829 ( .A(inst_register_registers[136]), .B(n3031), .C(
        inst_register_registers[40]), .D(n3032), .Y(n3033) );
  OAI21X1 U3830 ( .A(n3411), .B(n3561), .C(n3033), .Y(n3068) );
  NAND2X1 U3831 ( .A(instruction_ID[22]), .B(n4636), .Y(n3034) );
  NAND2X1 U3832 ( .A(instruction_ID[23]), .B(instruction_ID[22]), .Y(n3037) );
  NOR2X1 U3833 ( .A(n3035), .B(n3037), .Y(n3324) );
  AOI22X1 U3834 ( .A(inst_register_registers[72]), .B(n2806), .C(
        inst_register_registers[232]), .D(n3324), .Y(n3044) );
  NOR2X1 U3835 ( .A(n3036), .B(n3035), .Y(n3559) );
  AOI22X1 U3836 ( .A(inst_register_registers[104]), .B(n2808), .C(
        inst_register_registers[168]), .D(n3559), .Y(n3043) );
  NOR2X1 U3837 ( .A(n3040), .B(n3037), .Y(n3419) );
  NOR2X1 U3838 ( .A(n3040), .B(n3039), .Y(n3562) );
  AOI22X1 U3839 ( .A(inst_register_registers[200]), .B(n3038), .C(
        inst_register_registers[8]), .D(n3041), .Y(n3042) );
  NAND3X1 U3840 ( .A(n3044), .B(n3043), .C(n3042), .Y(n3067) );
  NOR2X1 U3841 ( .A(op_type_EX[0]), .B(n3045), .Y(n3063) );
  AOI22X1 U3842 ( .A(n3063), .B(read_register_2_EX[0]), .C(
        jump_inst_addr_EX[11]), .D(n3046), .Y(n3842) );
  AOI22X1 U3843 ( .A(n3063), .B(read_register_2_EX[2]), .C(
        jump_inst_addr_EX[13]), .D(n3046), .Y(n3840) );
  AOI22X1 U3844 ( .A(n3063), .B(read_register_2_EX[3]), .C(
        jump_inst_addr_EX[14]), .D(n3046), .Y(n3839) );
  AOI22X1 U3845 ( .A(n3063), .B(read_register_2_EX[4]), .C(n4414), .D(n3046), 
        .Y(n3838) );
  INVX1 U3846 ( .A(instruction_ID[17]), .Y(n4648) );
  AOI22X1 U3847 ( .A(n3063), .B(read_register_2_EX[1]), .C(
        jump_inst_addr_EX[12]), .D(n3046), .Y(n3841) );
  MUX2X1 U3848 ( .B(n4648), .A(instruction_ID[17]), .S(n3841), .Y(n3047) );
  OAI21X1 U3849 ( .A(instruction_ID[20]), .B(n3838), .C(n3047), .Y(n3048) );
  AOI21X1 U3850 ( .A(instruction_ID[20]), .B(n3838), .C(n3048), .Y(n3049) );
  OAI21X1 U3851 ( .A(instruction_ID[19]), .B(n3839), .C(n3049), .Y(n3050) );
  AOI21X1 U3852 ( .A(instruction_ID[19]), .B(n3839), .C(n3050), .Y(n3051) );
  OAI21X1 U3853 ( .A(instruction_ID[18]), .B(n3840), .C(n3051), .Y(n3052) );
  AOI21X1 U3854 ( .A(instruction_ID[18]), .B(n3840), .C(n3052), .Y(n3053) );
  OAI21X1 U3855 ( .A(instruction_ID[16]), .B(n3842), .C(n3053), .Y(n3054) );
  AOI21X1 U3856 ( .A(instruction_ID[16]), .B(n3842), .C(n3054), .Y(n3065) );
  MUX2X1 U3857 ( .B(n4638), .A(instruction_ID[22]), .S(n3841), .Y(n3055) );
  OAI21X1 U3858 ( .A(n3839), .B(instruction_ID[24]), .C(n3055), .Y(n3056) );
  AOI21X1 U3859 ( .A(n3839), .B(instruction_ID[24]), .C(n3056), .Y(n3057) );
  OAI21X1 U3860 ( .A(n3838), .B(instruction_ID[25]), .C(n3057), .Y(n3058) );
  AOI21X1 U3861 ( .A(n3838), .B(instruction_ID[25]), .C(n3058), .Y(n3059) );
  OAI21X1 U3862 ( .A(n3840), .B(instruction_ID[23]), .C(n3059), .Y(n3060) );
  AOI21X1 U3863 ( .A(n3840), .B(instruction_ID[23]), .C(n3060), .Y(n3061) );
  OAI21X1 U3864 ( .A(n3842), .B(instruction_ID[21]), .C(n3061), .Y(n3062) );
  AOI21X1 U3865 ( .A(n3842), .B(instruction_ID[21]), .C(n3062), .Y(n3064) );
  OAI21X1 U3866 ( .A(n3065), .B(n3064), .C(n3063), .Y(n3631) );
  AND2X2 U3867 ( .A(n3066), .B(n3631), .Y(n4705) );
  NAND2X1 U3868 ( .A(n4616), .B(n4705), .Y(n3933) );
  OAI21X1 U3869 ( .A(n3068), .B(n3067), .C(n2795), .Y(n3069) );
  AOI22X1 U3870 ( .A(inst_register_registers[66]), .B(n2806), .C(
        inst_register_registers[162]), .D(n3071), .Y(n3072) );
  OAI21X1 U3871 ( .A(n5129), .B(n3030), .C(n3072), .Y(n3078) );
  AOI22X1 U3872 ( .A(inst_register_registers[226]), .B(n3073), .C(
        inst_register_registers[2]), .D(n3041), .Y(n3076) );
  AOI22X1 U3873 ( .A(inst_register_registers[194]), .B(n3038), .C(
        inst_register_registers[130]), .D(n3564), .Y(n3075) );
  AOI22X1 U3874 ( .A(inst_register_registers[34]), .B(n3032), .C(
        inst_register_registers[98]), .D(n2808), .Y(n3074) );
  NAND3X1 U3875 ( .A(n3076), .B(n3075), .C(n3074), .Y(n3077) );
  OAI21X1 U3876 ( .A(n3078), .B(n3077), .C(n2795), .Y(n3079) );
  AOI22X1 U3877 ( .A(inst_register_registers[96]), .B(n2808), .C(
        inst_register_registers[192]), .D(n3038), .Y(n3081) );
  OAI21X1 U3878 ( .A(n3434), .B(n3030), .C(n3081), .Y(n3086) );
  AOI22X1 U3879 ( .A(inst_register_registers[128]), .B(n3031), .C(
        inst_register_registers[32]), .D(n3563), .Y(n3084) );
  AOI22X1 U3880 ( .A(inst_register_registers[160]), .B(n3071), .C(
        inst_register_registers[224]), .D(n3324), .Y(n3083) );
  AOI22X1 U3881 ( .A(inst_register_registers[64]), .B(n2806), .C(
        inst_register_registers[0]), .D(n3562), .Y(n3082) );
  NAND3X1 U3882 ( .A(n3084), .B(n3083), .C(n3082), .Y(n3085) );
  OAI21X1 U3883 ( .A(n3086), .B(n3085), .C(n2795), .Y(n3087) );
  AOI22X1 U3884 ( .A(inst_register_registers[235]), .B(n3073), .C(
        inst_register_registers[75]), .D(n2806), .Y(n3088) );
  OAI21X1 U3885 ( .A(n5156), .B(n3030), .C(n3088), .Y(n3093) );
  AOI22X1 U3886 ( .A(inst_register_registers[171]), .B(n3071), .C(
        inst_register_registers[43]), .D(n3563), .Y(n3091) );
  AOI22X1 U3887 ( .A(inst_register_registers[107]), .B(n2808), .C(
        inst_register_registers[203]), .D(n3038), .Y(n3090) );
  AOI22X1 U3888 ( .A(inst_register_registers[139]), .B(n3031), .C(
        inst_register_registers[11]), .D(n3562), .Y(n3089) );
  NAND3X1 U3889 ( .A(n3091), .B(n3090), .C(n3089), .Y(n3092) );
  OAI21X1 U3890 ( .A(n3093), .B(n3092), .C(n2795), .Y(n3094) );
  AOI22X1 U3891 ( .A(inst_register_registers[73]), .B(n2806), .C(
        inst_register_registers[9]), .D(n3041), .Y(n3095) );
  OAI21X1 U3892 ( .A(n5149), .B(n3561), .C(n3095), .Y(n3100) );
  AOI22X1 U3893 ( .A(inst_register_registers[105]), .B(n2808), .C(
        inst_register_registers[169]), .D(n3071), .Y(n3098) );
  AOI22X1 U3894 ( .A(inst_register_registers[233]), .B(n3073), .C(
        inst_register_registers[201]), .D(n3038), .Y(n3097) );
  AOI22X1 U3895 ( .A(inst_register_registers[41]), .B(n3032), .C(
        inst_register_registers[137]), .D(n3564), .Y(n3096) );
  NAND3X1 U3896 ( .A(n3098), .B(n3097), .C(n3096), .Y(n3099) );
  OAI21X1 U3897 ( .A(n3100), .B(n3099), .C(n2795), .Y(n3101) );
  AOI22X1 U3898 ( .A(inst_register_registers[37]), .B(n3032), .C(
        inst_register_registers[69]), .D(n2806), .Y(n3102) );
  OAI21X1 U3899 ( .A(n5138), .B(n3030), .C(n3102), .Y(n3107) );
  AOI22X1 U3900 ( .A(inst_register_registers[165]), .B(n3071), .C(
        inst_register_registers[101]), .D(n2808), .Y(n3105) );
  AOI22X1 U3901 ( .A(inst_register_registers[197]), .B(n3038), .C(
        inst_register_registers[229]), .D(n3073), .Y(n3104) );
  AOI22X1 U3902 ( .A(inst_register_registers[133]), .B(n3031), .C(
        inst_register_registers[5]), .D(n3562), .Y(n3103) );
  NAND3X1 U3903 ( .A(n3105), .B(n3104), .C(n3103), .Y(n3106) );
  OAI21X1 U3904 ( .A(n3107), .B(n3106), .C(n2795), .Y(n3108) );
  AOI22X1 U3905 ( .A(inst_register_registers[161]), .B(n3071), .C(
        inst_register_registers[1]), .D(n3041), .Y(n3109) );
  OAI21X1 U3906 ( .A(n5126), .B(n3030), .C(n3109), .Y(n3114) );
  AOI22X1 U3907 ( .A(inst_register_registers[97]), .B(n2808), .C(
        inst_register_registers[193]), .D(n3038), .Y(n3112) );
  AOI22X1 U3908 ( .A(inst_register_registers[225]), .B(n3073), .C(
        inst_register_registers[65]), .D(n2806), .Y(n3111) );
  AOI22X1 U3909 ( .A(inst_register_registers[129]), .B(n3031), .C(
        inst_register_registers[33]), .D(n3563), .Y(n3110) );
  NAND3X1 U3910 ( .A(n3112), .B(n3111), .C(n3110), .Y(n3113) );
  OAI21X1 U3911 ( .A(n3114), .B(n3113), .C(n2795), .Y(n3115) );
  AOI22X1 U3912 ( .A(inst_register_registers[7]), .B(n3041), .C(
        inst_register_registers[231]), .D(n3324), .Y(n3116) );
  OAI21X1 U3913 ( .A(n5144), .B(n3030), .C(n3116), .Y(n3121) );
  AOI22X1 U3914 ( .A(inst_register_registers[167]), .B(n3071), .C(
        inst_register_registers[39]), .D(n3032), .Y(n3119) );
  AOI22X1 U3915 ( .A(inst_register_registers[199]), .B(n3038), .C(
        inst_register_registers[71]), .D(n2806), .Y(n3118) );
  AOI22X1 U3916 ( .A(inst_register_registers[135]), .B(n3031), .C(
        inst_register_registers[103]), .D(n2808), .Y(n3117) );
  NAND3X1 U3917 ( .A(n3119), .B(n3118), .C(n3117), .Y(n3120) );
  OAI21X1 U3918 ( .A(n3121), .B(n3120), .C(n2795), .Y(n3122) );
  AOI22X1 U3919 ( .A(inst_register_registers[230]), .B(n3073), .C(
        inst_register_registers[38]), .D(n3563), .Y(n3123) );
  OAI21X1 U3920 ( .A(n5141), .B(n3030), .C(n3123), .Y(n3128) );
  AOI22X1 U3921 ( .A(inst_register_registers[6]), .B(n3041), .C(
        inst_register_registers[198]), .D(n3038), .Y(n3126) );
  AOI22X1 U3922 ( .A(inst_register_registers[134]), .B(n3031), .C(
        inst_register_registers[102]), .D(n2808), .Y(n3125) );
  AOI22X1 U3923 ( .A(inst_register_registers[166]), .B(n3071), .C(
        inst_register_registers[70]), .D(n2806), .Y(n3124) );
  NAND3X1 U3924 ( .A(n3126), .B(n3125), .C(n3124), .Y(n3127) );
  OAI21X1 U3925 ( .A(n3128), .B(n3127), .C(n2795), .Y(n3129) );
  AOI22X1 U3926 ( .A(inst_register_registers[172]), .B(n3071), .C(
        inst_register_registers[44]), .D(n3032), .Y(n3130) );
  OAI21X1 U3927 ( .A(n5159), .B(n3030), .C(n3130), .Y(n3135) );
  AOI22X1 U3928 ( .A(inst_register_registers[12]), .B(n3041), .C(
        inst_register_registers[236]), .D(n3073), .Y(n3133) );
  AOI22X1 U3929 ( .A(inst_register_registers[140]), .B(n3031), .C(
        inst_register_registers[204]), .D(n3419), .Y(n3132) );
  AOI22X1 U3930 ( .A(inst_register_registers[108]), .B(n2808), .C(
        inst_register_registers[76]), .D(n2806), .Y(n3131) );
  NAND3X1 U3931 ( .A(n3133), .B(n3132), .C(n3131), .Y(n3134) );
  OAI21X1 U3932 ( .A(n3135), .B(n3134), .C(n2795), .Y(n3136) );
  MUX2X1 U3933 ( .B(alu_result_WB[31]), .A(mem_read_data_WB[31]), .S(n3534), 
        .Y(n3949) );
  INVX1 U3934 ( .A(instruction_ID[18]), .Y(n4646) );
  INVX1 U3935 ( .A(instruction_ID[20]), .Y(n4642) );
  AOI22X1 U3936 ( .A(reg_write_address_WB[4]), .B(instruction_ID[20]), .C(
        n4642), .D(n3137), .Y(n3144) );
  AOI22X1 U3937 ( .A(reg_write_address_WB[1]), .B(n4648), .C(
        instruction_ID[17]), .D(n5428), .Y(n3138) );
  OAI21X1 U3938 ( .A(instruction_ID[19]), .B(n3139), .C(n3138), .Y(n3141) );
  INVX1 U3939 ( .A(instruction_ID[19]), .Y(n4644) );
  OAI21X1 U3940 ( .A(reg_write_address_WB[3]), .B(n4644), .C(n5202), .Y(n3140)
         );
  NOR2X1 U3941 ( .A(n3141), .B(n3140), .Y(n3142) );
  OAI21X1 U3942 ( .A(instruction_ID[18]), .B(n5391), .C(n3142), .Y(n3143) );
  NOR2X1 U3943 ( .A(n3144), .B(n3143), .Y(n3145) );
  OAI21X1 U3944 ( .A(reg_write_address_WB[2]), .B(n4646), .C(n3145), .Y(n3146)
         );
  AOI21X1 U3945 ( .A(n5201), .B(instruction_ID[16]), .C(n3146), .Y(n3147) );
  OAI21X1 U3946 ( .A(n5201), .B(instruction_ID[16]), .C(n3147), .Y(n3537) );
  INVX1 U3947 ( .A(instruction_ID[16]), .Y(n4650) );
  NAND2X1 U3948 ( .A(n4650), .B(n3148), .Y(n3153) );
  NAND2X1 U3949 ( .A(instruction_ID[18]), .B(n4648), .Y(n3149) );
  NAND2X1 U3950 ( .A(instruction_ID[16]), .B(n3148), .Y(n3155) );
  AOI22X1 U3951 ( .A(n2802), .B(inst_register_registers[159]), .C(n2801), .D(
        inst_register_registers[191]), .Y(n3150) );
  OAI21X1 U3952 ( .A(n3949), .B(n3537), .C(n3150), .Y(n3161) );
  NAND2X1 U3953 ( .A(n4646), .B(n4648), .Y(n3151) );
  AOI22X1 U3954 ( .A(n2803), .B(inst_register_registers[31]), .C(n2804), .D(
        inst_register_registers[63]), .Y(n3159) );
  NAND2X1 U3955 ( .A(instruction_ID[17]), .B(n4646), .Y(n3152) );
  NOR2X1 U3956 ( .A(n3152), .B(n3155), .Y(n3535) );
  AOI22X1 U3957 ( .A(n2805), .B(inst_register_registers[95]), .C(n3535), .D(
        inst_register_registers[127]), .Y(n3158) );
  NAND2X1 U3958 ( .A(instruction_ID[18]), .B(instruction_ID[17]), .Y(n3154) );
  NOR2X1 U3959 ( .A(n3155), .B(n3154), .Y(n3552) );
  AOI22X1 U3960 ( .A(n2807), .B(inst_register_registers[223]), .C(n3156), .D(
        inst_register_registers[255]), .Y(n3157) );
  NAND3X1 U3961 ( .A(n3159), .B(n3158), .C(n3157), .Y(n3160) );
  OAI21X1 U3962 ( .A(n3161), .B(n3160), .C(n2795), .Y(n3162) );
  AOI22X1 U3963 ( .A(inst_register_registers[31]), .B(n3041), .C(
        inst_register_registers[95]), .D(n2806), .Y(n3163) );
  OAI21X1 U3964 ( .A(n3949), .B(n3030), .C(n3163), .Y(n3168) );
  AOI22X1 U3965 ( .A(inst_register_registers[127]), .B(n2808), .C(
        inst_register_registers[255]), .D(n3324), .Y(n3166) );
  AOI22X1 U3966 ( .A(inst_register_registers[63]), .B(n3032), .C(
        inst_register_registers[223]), .D(n3419), .Y(n3165) );
  AOI22X1 U3967 ( .A(inst_register_registers[191]), .B(n3071), .C(
        inst_register_registers[159]), .D(n3564), .Y(n3164) );
  NAND3X1 U3968 ( .A(n3166), .B(n3165), .C(n3164), .Y(n3167) );
  OAI21X1 U3969 ( .A(n3168), .B(n3167), .C(n2795), .Y(n3169) );
  AOI22X1 U3970 ( .A(inst_register_registers[170]), .B(n3071), .C(
        inst_register_registers[202]), .D(n3038), .Y(n3170) );
  OAI21X1 U3971 ( .A(n5152), .B(n3561), .C(n3170), .Y(n3175) );
  AOI22X1 U3972 ( .A(inst_register_registers[234]), .B(n3073), .C(
        inst_register_registers[42]), .D(n3563), .Y(n3173) );
  AOI22X1 U3973 ( .A(inst_register_registers[138]), .B(n3031), .C(
        inst_register_registers[106]), .D(n2808), .Y(n3172) );
  AOI22X1 U3974 ( .A(inst_register_registers[10]), .B(n3041), .C(
        inst_register_registers[74]), .D(n2806), .Y(n3171) );
  NAND3X1 U3975 ( .A(n3173), .B(n3172), .C(n3171), .Y(n3174) );
  OAI21X1 U3976 ( .A(n3175), .B(n3174), .C(n2795), .Y(n3176) );
  AOI22X1 U3977 ( .A(inst_register_registers[227]), .B(n3073), .C(
        inst_register_registers[67]), .D(n2806), .Y(n3177) );
  OAI21X1 U3978 ( .A(n5132), .B(n3030), .C(n3177), .Y(n3182) );
  AOI22X1 U3979 ( .A(inst_register_registers[99]), .B(n2808), .C(
        inst_register_registers[35]), .D(n3563), .Y(n3180) );
  AOI22X1 U3980 ( .A(inst_register_registers[3]), .B(n3041), .C(
        inst_register_registers[195]), .D(n3038), .Y(n3179) );
  AOI22X1 U3981 ( .A(inst_register_registers[163]), .B(n3071), .C(
        inst_register_registers[131]), .D(n3564), .Y(n3178) );
  NAND3X1 U3982 ( .A(n3180), .B(n3179), .C(n3178), .Y(n3181) );
  OAI21X1 U3983 ( .A(n3182), .B(n3181), .C(n2795), .Y(n3183) );
  AOI22X1 U3984 ( .A(inst_register_registers[36]), .B(n3032), .C(
        inst_register_registers[228]), .D(n3324), .Y(n3184) );
  OAI21X1 U3985 ( .A(n5135), .B(n3030), .C(n3184), .Y(n3189) );
  AOI22X1 U3986 ( .A(inst_register_registers[100]), .B(n2808), .C(
        inst_register_registers[196]), .D(n3038), .Y(n3187) );
  AOI22X1 U3987 ( .A(inst_register_registers[68]), .B(n2806), .C(
        inst_register_registers[132]), .D(n3564), .Y(n3186) );
  AOI22X1 U3988 ( .A(inst_register_registers[164]), .B(n3071), .C(
        inst_register_registers[4]), .D(n3041), .Y(n3185) );
  NAND3X1 U3989 ( .A(n3187), .B(n3186), .C(n3185), .Y(n3188) );
  OAI21X1 U3990 ( .A(n3189), .B(n3188), .C(n2795), .Y(n3190) );
  FAX1 U3991 ( .A(n4071), .B(n3192), .C(n3191), .YC(n4026), .YS(n3196) );
  NAND2X1 U3992 ( .A(n4071), .B(n4083), .Y(n3194) );
  OAI21X1 U3993 ( .A(n4083), .B(n4071), .C(n3739), .Y(n3193) );
  OAI21X1 U3994 ( .A(n3194), .B(n4047), .C(n3193), .Y(n3195) );
  AOI21X1 U3995 ( .A(n4263), .B(n3196), .C(n3195), .Y(n3197) );
  FAX1 U3996 ( .A(n4072), .B(n3199), .C(n3198), .YC(n3191), .YS(n3203) );
  NAND2X1 U3997 ( .A(n4072), .B(n4077), .Y(n3201) );
  OAI21X1 U3998 ( .A(n4077), .B(n4072), .C(n3739), .Y(n3200) );
  OAI21X1 U3999 ( .A(n3201), .B(n4047), .C(n3200), .Y(n3202) );
  AOI21X1 U4000 ( .A(n4263), .B(n3203), .C(n3202), .Y(n3204) );
  MUX2X1 U4001 ( .B(alu_result_WB[22]), .A(mem_read_data_WB[22]), .S(n3534), 
        .Y(n3685) );
  AOI22X1 U4002 ( .A(n2802), .B(inst_register_registers[150]), .C(n2801), .D(
        inst_register_registers[182]), .Y(n3206) );
  OAI21X1 U4003 ( .A(n3685), .B(n3148), .C(n3206), .Y(n3214) );
  AOI22X1 U4004 ( .A(n3207), .B(inst_register_registers[118]), .C(n3552), .D(
        inst_register_registers[246]), .Y(n3212) );
  AOI22X1 U4005 ( .A(n2805), .B(inst_register_registers[86]), .C(n2803), .D(
        inst_register_registers[22]), .Y(n3211) );
  AOI22X1 U4006 ( .A(n2807), .B(inst_register_registers[214]), .C(n2804), .D(
        inst_register_registers[54]), .Y(n3210) );
  NAND3X1 U4007 ( .A(n3212), .B(n3211), .C(n3210), .Y(n3213) );
  OAI21X1 U4008 ( .A(n3214), .B(n3213), .C(n2795), .Y(n3215) );
  MUX2X1 U4009 ( .B(alu_result_WB[23]), .A(mem_read_data_WB[23]), .S(n3534), 
        .Y(n3696) );
  AOI22X1 U4010 ( .A(inst_register_registers[87]), .B(n2806), .C(
        inst_register_registers[247]), .D(n3324), .Y(n3216) );
  OAI21X1 U4011 ( .A(n3696), .B(n3030), .C(n3216), .Y(n3221) );
  AOI22X1 U4012 ( .A(inst_register_registers[55]), .B(n3032), .C(
        inst_register_registers[151]), .D(n3031), .Y(n3219) );
  AOI22X1 U4013 ( .A(inst_register_registers[23]), .B(n3041), .C(
        inst_register_registers[119]), .D(n2808), .Y(n3218) );
  AOI22X1 U4014 ( .A(inst_register_registers[183]), .B(n3071), .C(
        inst_register_registers[215]), .D(n3419), .Y(n3217) );
  NAND3X1 U4015 ( .A(n3219), .B(n3218), .C(n3217), .Y(n3220) );
  OAI21X1 U4016 ( .A(n3221), .B(n3220), .C(n2795), .Y(n3222) );
  MUX2X1 U4017 ( .B(alu_result_WB[21]), .A(mem_read_data_WB[21]), .S(n3534), 
        .Y(n3670) );
  AOI22X1 U4018 ( .A(n2804), .B(inst_register_registers[53]), .C(n2801), .D(
        inst_register_registers[181]), .Y(n3224) );
  OAI21X1 U4019 ( .A(n3670), .B(n3148), .C(n3224), .Y(n3229) );
  AOI22X1 U4020 ( .A(n3207), .B(inst_register_registers[117]), .C(n2802), .D(
        inst_register_registers[149]), .Y(n3227) );
  AOI22X1 U4021 ( .A(n2805), .B(inst_register_registers[85]), .C(n2803), .D(
        inst_register_registers[21]), .Y(n3226) );
  AOI22X1 U4022 ( .A(n2807), .B(inst_register_registers[213]), .C(n3156), .D(
        inst_register_registers[245]), .Y(n3225) );
  NAND3X1 U4023 ( .A(n3227), .B(n3226), .C(n3225), .Y(n3228) );
  OAI21X1 U4024 ( .A(n3229), .B(n3228), .C(n2795), .Y(n3230) );
  MUX2X1 U4025 ( .B(alu_result_WB[25]), .A(mem_read_data_WB[25]), .S(n3534), 
        .Y(n5189) );
  AOI22X1 U4026 ( .A(inst_register_registers[185]), .B(n3559), .C(
        inst_register_registers[121]), .D(n2808), .Y(n3231) );
  OAI21X1 U4027 ( .A(n5189), .B(n3030), .C(n3231), .Y(n3236) );
  AOI22X1 U4028 ( .A(inst_register_registers[217]), .B(n3038), .C(
        inst_register_registers[57]), .D(n3032), .Y(n3234) );
  AOI22X1 U4029 ( .A(inst_register_registers[153]), .B(n3031), .C(
        inst_register_registers[89]), .D(n2806), .Y(n3233) );
  AOI22X1 U4030 ( .A(inst_register_registers[25]), .B(n3041), .C(
        inst_register_registers[249]), .D(n3324), .Y(n3232) );
  NAND3X1 U4031 ( .A(n3234), .B(n3233), .C(n3232), .Y(n3235) );
  OAI21X1 U4032 ( .A(n3236), .B(n3235), .C(n2795), .Y(n3237) );
  MUX2X1 U4033 ( .B(alu_result_WB[20]), .A(mem_read_data_WB[20]), .S(n3534), 
        .Y(n3674) );
  AOI22X1 U4034 ( .A(n2805), .B(inst_register_registers[84]), .C(n3156), .D(
        inst_register_registers[244]), .Y(n3238) );
  OAI21X1 U4035 ( .A(n3674), .B(n3148), .C(n3238), .Y(n3243) );
  AOI22X1 U4036 ( .A(n2807), .B(inst_register_registers[212]), .C(n2802), .D(
        inst_register_registers[148]), .Y(n3241) );
  AOI22X1 U4037 ( .A(n2803), .B(inst_register_registers[20]), .C(n2801), .D(
        inst_register_registers[180]), .Y(n3240) );
  AOI22X1 U4038 ( .A(n3207), .B(inst_register_registers[116]), .C(n2804), .D(
        inst_register_registers[52]), .Y(n3239) );
  NAND3X1 U4039 ( .A(n3241), .B(n3240), .C(n3239), .Y(n3242) );
  OAI21X1 U4040 ( .A(n3243), .B(n3242), .C(n2795), .Y(n3244) );
  MUX2X1 U4041 ( .B(alu_result_WB[24]), .A(mem_read_data_WB[24]), .S(n3534), 
        .Y(n5186) );
  AOI22X1 U4042 ( .A(n2805), .B(inst_register_registers[88]), .C(n2807), .D(
        inst_register_registers[216]), .Y(n3246) );
  OAI21X1 U4043 ( .A(n5186), .B(n3148), .C(n3246), .Y(n3251) );
  AOI22X1 U4044 ( .A(n2801), .B(inst_register_registers[184]), .C(n3552), .D(
        inst_register_registers[248]), .Y(n3249) );
  AOI22X1 U4045 ( .A(n3207), .B(inst_register_registers[120]), .C(n2802), .D(
        inst_register_registers[152]), .Y(n3248) );
  AOI22X1 U4046 ( .A(n2803), .B(inst_register_registers[24]), .C(n2804), .D(
        inst_register_registers[56]), .Y(n3247) );
  NAND3X1 U4047 ( .A(n3249), .B(n3248), .C(n3247), .Y(n3250) );
  OAI21X1 U4048 ( .A(n3251), .B(n3250), .C(n2795), .Y(n3252) );
  AOI22X1 U4049 ( .A(inst_register_registers[118]), .B(n2808), .C(
        inst_register_registers[22]), .D(n3041), .Y(n3253) );
  OAI21X1 U4050 ( .A(n3685), .B(n3030), .C(n3253), .Y(n3258) );
  AOI22X1 U4051 ( .A(inst_register_registers[86]), .B(n2806), .C(
        inst_register_registers[182]), .D(n3559), .Y(n3256) );
  AOI22X1 U4052 ( .A(inst_register_registers[214]), .B(n3038), .C(
        inst_register_registers[150]), .D(n3564), .Y(n3255) );
  AOI22X1 U4053 ( .A(inst_register_registers[246]), .B(n3073), .C(
        inst_register_registers[54]), .D(n3032), .Y(n3254) );
  NAND3X1 U4054 ( .A(n3256), .B(n3255), .C(n3254), .Y(n3257) );
  OAI21X1 U4055 ( .A(n3258), .B(n3257), .C(n2795), .Y(n3259) );
  AOI22X1 U4056 ( .A(inst_register_registers[184]), .B(n3071), .C(
        inst_register_registers[24]), .D(n3562), .Y(n3260) );
  OAI21X1 U4057 ( .A(n5186), .B(n3030), .C(n3260), .Y(n3265) );
  AOI22X1 U4058 ( .A(inst_register_registers[120]), .B(n2808), .C(
        inst_register_registers[216]), .D(n3419), .Y(n3263) );
  AOI22X1 U4059 ( .A(inst_register_registers[152]), .B(n3031), .C(
        inst_register_registers[56]), .D(n3032), .Y(n3262) );
  AOI22X1 U4060 ( .A(inst_register_registers[248]), .B(n3073), .C(
        inst_register_registers[88]), .D(n2806), .Y(n3261) );
  NAND3X1 U4061 ( .A(n3263), .B(n3262), .C(n3261), .Y(n3264) );
  OAI21X1 U4062 ( .A(n3265), .B(n3264), .C(n2795), .Y(n3266) );
  AOI22X1 U4063 ( .A(inst_register_registers[20]), .B(n3041), .C(
        inst_register_registers[52]), .D(n3032), .Y(n3267) );
  OAI21X1 U4064 ( .A(n3674), .B(n3030), .C(n3267), .Y(n3272) );
  AOI22X1 U4065 ( .A(inst_register_registers[212]), .B(n3038), .C(
        inst_register_registers[148]), .D(n3031), .Y(n3270) );
  AOI22X1 U4066 ( .A(inst_register_registers[116]), .B(n2808), .C(
        inst_register_registers[244]), .D(n3324), .Y(n3269) );
  AOI22X1 U4067 ( .A(inst_register_registers[180]), .B(n3071), .C(
        inst_register_registers[84]), .D(n2806), .Y(n3268) );
  NAND3X1 U4068 ( .A(n3270), .B(n3269), .C(n3268), .Y(n3271) );
  OAI21X1 U4069 ( .A(n3272), .B(n3271), .C(n2795), .Y(n3273) );
  AOI22X1 U4070 ( .A(n2807), .B(inst_register_registers[215]), .C(n3552), .D(
        inst_register_registers[247]), .Y(n3274) );
  OAI21X1 U4071 ( .A(n3696), .B(n3148), .C(n3274), .Y(n3279) );
  AOI22X1 U4072 ( .A(n2803), .B(inst_register_registers[23]), .C(n2804), .D(
        inst_register_registers[55]), .Y(n3277) );
  AOI22X1 U4073 ( .A(n2805), .B(inst_register_registers[87]), .C(n2802), .D(
        inst_register_registers[151]), .Y(n3276) );
  AOI22X1 U4074 ( .A(n3207), .B(inst_register_registers[119]), .C(n2801), .D(
        inst_register_registers[183]), .Y(n3275) );
  NAND3X1 U4075 ( .A(n3277), .B(n3276), .C(n3275), .Y(n3278) );
  OAI21X1 U4076 ( .A(n3279), .B(n3278), .C(n2795), .Y(n3280) );
  AOI22X1 U4077 ( .A(inst_register_registers[110]), .B(n2808), .C(
        inst_register_registers[206]), .D(n3038), .Y(n3281) );
  OAI21X1 U4078 ( .A(n3442), .B(n3561), .C(n3281), .Y(n3286) );
  AOI22X1 U4079 ( .A(inst_register_registers[174]), .B(n3071), .C(
        inst_register_registers[238]), .D(n3324), .Y(n3284) );
  AOI22X1 U4080 ( .A(inst_register_registers[78]), .B(n2806), .C(
        inst_register_registers[14]), .D(n3562), .Y(n3283) );
  AOI22X1 U4081 ( .A(inst_register_registers[142]), .B(n3031), .C(
        inst_register_registers[46]), .D(n3032), .Y(n3282) );
  NAND3X1 U4082 ( .A(n3284), .B(n3283), .C(n3282), .Y(n3285) );
  OAI21X1 U4083 ( .A(n3286), .B(n3285), .C(n2795), .Y(n3287) );
  AOI22X1 U4084 ( .A(inst_register_registers[173]), .B(n3071), .C(
        inst_register_registers[205]), .D(n3419), .Y(n3288) );
  OAI21X1 U4085 ( .A(n5162), .B(n3030), .C(n3288), .Y(n3293) );
  AOI22X1 U4086 ( .A(inst_register_registers[141]), .B(n3031), .C(
        inst_register_registers[45]), .D(n3563), .Y(n3291) );
  AOI22X1 U4087 ( .A(inst_register_registers[77]), .B(n2806), .C(
        inst_register_registers[13]), .D(n3562), .Y(n3290) );
  AOI22X1 U4088 ( .A(inst_register_registers[237]), .B(n3073), .C(
        inst_register_registers[109]), .D(n2808), .Y(n3289) );
  NAND3X1 U4089 ( .A(n3291), .B(n3290), .C(n3289), .Y(n3292) );
  OAI21X1 U4090 ( .A(n3293), .B(n3292), .C(n2795), .Y(n3294) );
  MUX2X1 U4091 ( .B(alu_result_WB[19]), .A(mem_read_data_WB[19]), .S(n3534), 
        .Y(n3652) );
  AOI22X1 U4092 ( .A(inst_register_registers[19]), .B(n3041), .C(
        inst_register_registers[83]), .D(n2806), .Y(n3295) );
  OAI21X1 U4093 ( .A(n3652), .B(n3561), .C(n3295), .Y(n3300) );
  AOI22X1 U4094 ( .A(inst_register_registers[51]), .B(n3032), .C(
        inst_register_registers[179]), .D(n3559), .Y(n3298) );
  AOI22X1 U4095 ( .A(inst_register_registers[243]), .B(n3073), .C(
        inst_register_registers[115]), .D(n2808), .Y(n3297) );
  AOI22X1 U4096 ( .A(inst_register_registers[211]), .B(n3038), .C(
        inst_register_registers[147]), .D(n3564), .Y(n3296) );
  NAND3X1 U4097 ( .A(n3298), .B(n3297), .C(n3296), .Y(n3299) );
  OAI21X1 U4098 ( .A(n3300), .B(n3299), .C(n2795), .Y(n3301) );
  MUX2X1 U4099 ( .B(alu_result_WB[26]), .A(mem_read_data_WB[26]), .S(n3534), 
        .Y(n5192) );
  AOI22X1 U4100 ( .A(n3535), .B(inst_register_registers[122]), .C(n2801), .D(
        inst_register_registers[186]), .Y(n3302) );
  OAI21X1 U4101 ( .A(n5192), .B(n3148), .C(n3302), .Y(n3307) );
  AOI22X1 U4102 ( .A(n2805), .B(inst_register_registers[90]), .C(n2802), .D(
        inst_register_registers[154]), .Y(n3305) );
  AOI22X1 U4103 ( .A(n2807), .B(inst_register_registers[218]), .C(n3156), .D(
        inst_register_registers[250]), .Y(n3304) );
  AOI22X1 U4104 ( .A(n2803), .B(inst_register_registers[26]), .C(n2804), .D(
        inst_register_registers[58]), .Y(n3303) );
  NAND3X1 U4105 ( .A(n3305), .B(n3304), .C(n3303), .Y(n3306) );
  OAI21X1 U4106 ( .A(n3307), .B(n3306), .C(n2795), .Y(n3308) );
  AOI22X1 U4107 ( .A(n2807), .B(inst_register_registers[217]), .C(n2804), .D(
        inst_register_registers[57]), .Y(n3309) );
  OAI21X1 U4108 ( .A(n5189), .B(n3148), .C(n3309), .Y(n3314) );
  AOI22X1 U4109 ( .A(n2803), .B(inst_register_registers[25]), .C(n2802), .D(
        inst_register_registers[153]), .Y(n3312) );
  AOI22X1 U4110 ( .A(n2801), .B(inst_register_registers[185]), .C(n3156), .D(
        inst_register_registers[249]), .Y(n3311) );
  AOI22X1 U4111 ( .A(n2805), .B(inst_register_registers[89]), .C(n3535), .D(
        inst_register_registers[121]), .Y(n3310) );
  NAND3X1 U4112 ( .A(n3312), .B(n3311), .C(n3310), .Y(n3313) );
  OAI21X1 U4113 ( .A(n3314), .B(n3313), .C(n2795), .Y(n3315) );
  AOI22X1 U4114 ( .A(inst_register_registers[218]), .B(n3038), .C(
        inst_register_registers[58]), .D(n3032), .Y(n3316) );
  OAI21X1 U4115 ( .A(n5192), .B(n3030), .C(n3316), .Y(n3321) );
  AOI22X1 U4116 ( .A(inst_register_registers[250]), .B(n3073), .C(
        inst_register_registers[26]), .D(n3041), .Y(n3319) );
  AOI22X1 U4117 ( .A(inst_register_registers[186]), .B(n3071), .C(
        inst_register_registers[122]), .D(n2808), .Y(n3318) );
  AOI22X1 U4118 ( .A(inst_register_registers[154]), .B(n3031), .C(
        inst_register_registers[90]), .D(n2806), .Y(n3317) );
  NAND3X1 U4119 ( .A(n3319), .B(n3318), .C(n3317), .Y(n3320) );
  OAI21X1 U4120 ( .A(n3321), .B(n3320), .C(n2795), .Y(n3322) );
  AOI22X1 U4121 ( .A(inst_register_registers[85]), .B(n2806), .C(
        inst_register_registers[53]), .D(n3032), .Y(n3323) );
  OAI21X1 U4122 ( .A(n3670), .B(n3030), .C(n3323), .Y(n3329) );
  AOI22X1 U4123 ( .A(inst_register_registers[21]), .B(n3041), .C(
        inst_register_registers[245]), .D(n3324), .Y(n3327) );
  AOI22X1 U4124 ( .A(inst_register_registers[213]), .B(n3038), .C(
        inst_register_registers[181]), .D(n3559), .Y(n3326) );
  AOI22X1 U4125 ( .A(inst_register_registers[117]), .B(n2808), .C(
        inst_register_registers[149]), .D(n3564), .Y(n3325) );
  NAND3X1 U4126 ( .A(n3327), .B(n3326), .C(n3325), .Y(n3328) );
  OAI21X1 U4127 ( .A(n3329), .B(n3328), .C(n2795), .Y(n3330) );
  MUX2X1 U4128 ( .B(alu_result_WB[27]), .A(mem_read_data_WB[27]), .S(n3534), 
        .Y(n5195) );
  AOI22X1 U4129 ( .A(inst_register_registers[251]), .B(n3073), .C(
        inst_register_registers[27]), .D(n3041), .Y(n3331) );
  OAI21X1 U4130 ( .A(n5195), .B(n3561), .C(n3331), .Y(n3336) );
  AOI22X1 U4131 ( .A(inst_register_registers[155]), .B(n3031), .C(
        inst_register_registers[187]), .D(n3071), .Y(n3334) );
  AOI22X1 U4132 ( .A(inst_register_registers[59]), .B(n3032), .C(
        inst_register_registers[91]), .D(n2806), .Y(n3333) );
  AOI22X1 U4133 ( .A(inst_register_registers[123]), .B(n2808), .C(
        inst_register_registers[219]), .D(n3419), .Y(n3332) );
  NAND3X1 U4134 ( .A(n3334), .B(n3333), .C(n3332), .Y(n3335) );
  OAI21X1 U4135 ( .A(n3336), .B(n3335), .C(n2795), .Y(n3337) );
  MUX2X1 U4136 ( .B(alu_result_WB[28]), .A(mem_read_data_WB[28]), .S(n3534), 
        .Y(n5198) );
  AOI22X1 U4137 ( .A(n2807), .B(inst_register_registers[220]), .C(n2802), .D(
        inst_register_registers[156]), .Y(n3338) );
  OAI21X1 U4138 ( .A(n5198), .B(n3537), .C(n3338), .Y(n3343) );
  AOI22X1 U4139 ( .A(n2803), .B(inst_register_registers[28]), .C(n3535), .D(
        inst_register_registers[124]), .Y(n3341) );
  AOI22X1 U4140 ( .A(n2801), .B(inst_register_registers[188]), .C(n3156), .D(
        inst_register_registers[252]), .Y(n3340) );
  AOI22X1 U4141 ( .A(n2805), .B(inst_register_registers[92]), .C(n2804), .D(
        inst_register_registers[60]), .Y(n3339) );
  NAND3X1 U4142 ( .A(n3341), .B(n3340), .C(n3339), .Y(n3342) );
  OAI21X1 U4143 ( .A(n3343), .B(n3342), .C(n2795), .Y(n3344) );
  AOI22X1 U4144 ( .A(inst_register_registers[112]), .B(n2808), .C(
        inst_register_registers[144]), .D(n3031), .Y(n3345) );
  OAI21X1 U4145 ( .A(n3506), .B(n3561), .C(n3345), .Y(n3350) );
  AOI22X1 U4146 ( .A(inst_register_registers[240]), .B(n3073), .C(
        inst_register_registers[208]), .D(n3419), .Y(n3348) );
  AOI22X1 U4147 ( .A(inst_register_registers[176]), .B(n3071), .C(
        inst_register_registers[80]), .D(n2806), .Y(n3347) );
  AOI22X1 U4148 ( .A(inst_register_registers[48]), .B(n3032), .C(
        inst_register_registers[16]), .D(n3562), .Y(n3346) );
  NAND3X1 U4149 ( .A(n3348), .B(n3347), .C(n3346), .Y(n3349) );
  OAI21X1 U4150 ( .A(n3350), .B(n3349), .C(n2795), .Y(n3351) );
  MUX2X1 U4151 ( .B(alu_result_WB[17]), .A(mem_read_data_WB[17]), .S(n3534), 
        .Y(n5171) );
  AOI22X1 U4152 ( .A(inst_register_registers[113]), .B(n2808), .C(
        inst_register_registers[49]), .D(n3032), .Y(n3352) );
  OAI21X1 U4153 ( .A(n5171), .B(n3030), .C(n3352), .Y(n3357) );
  AOI22X1 U4154 ( .A(inst_register_registers[81]), .B(n2806), .C(
        inst_register_registers[145]), .D(n3031), .Y(n3355) );
  AOI22X1 U4155 ( .A(inst_register_registers[17]), .B(n3041), .C(
        inst_register_registers[177]), .D(n3559), .Y(n3354) );
  AOI22X1 U4156 ( .A(inst_register_registers[241]), .B(n3073), .C(
        inst_register_registers[209]), .D(n3419), .Y(n3353) );
  NAND3X1 U4157 ( .A(n3355), .B(n3354), .C(n3353), .Y(n3356) );
  OAI21X1 U4158 ( .A(n3357), .B(n3356), .C(n2795), .Y(n3358) );
  AOI22X1 U4159 ( .A(inst_register_registers[143]), .B(n3031), .C(
        inst_register_registers[239]), .D(n3073), .Y(n3359) );
  OAI21X1 U4160 ( .A(n3389), .B(n3561), .C(n3359), .Y(n3364) );
  AOI22X1 U4161 ( .A(inst_register_registers[79]), .B(n2806), .C(
        inst_register_registers[207]), .D(n3419), .Y(n3362) );
  AOI22X1 U4162 ( .A(inst_register_registers[47]), .B(n3032), .C(
        inst_register_registers[175]), .D(n3559), .Y(n3361) );
  AOI22X1 U4163 ( .A(inst_register_registers[111]), .B(n2808), .C(
        inst_register_registers[15]), .D(n3562), .Y(n3360) );
  NAND3X1 U4164 ( .A(n3362), .B(n3361), .C(n3360), .Y(n3363) );
  OAI21X1 U4165 ( .A(n3364), .B(n3363), .C(n2795), .Y(n3365) );
  AOI22X1 U4166 ( .A(n2805), .B(inst_register_registers[91]), .C(n2807), .D(
        inst_register_registers[219]), .Y(n3366) );
  OAI21X1 U4167 ( .A(n5195), .B(n3537), .C(n3366), .Y(n3371) );
  AOI22X1 U4168 ( .A(n2802), .B(inst_register_registers[155]), .C(n3156), .D(
        inst_register_registers[251]), .Y(n3369) );
  AOI22X1 U4169 ( .A(n2803), .B(inst_register_registers[27]), .C(n3535), .D(
        inst_register_registers[123]), .Y(n3368) );
  AOI22X1 U4170 ( .A(n2804), .B(inst_register_registers[59]), .C(n2801), .D(
        inst_register_registers[187]), .Y(n3367) );
  NAND3X1 U4171 ( .A(n3369), .B(n3368), .C(n3367), .Y(n3370) );
  OAI21X1 U4172 ( .A(n3371), .B(n3370), .C(n2795), .Y(n3372) );
  MUX2X1 U4173 ( .B(alu_result_WB[18]), .A(mem_read_data_WB[18]), .S(n3534), 
        .Y(n3656) );
  AOI22X1 U4174 ( .A(inst_register_registers[82]), .B(n2806), .C(
        inst_register_registers[242]), .D(n3073), .Y(n3373) );
  OAI21X1 U4175 ( .A(n3656), .B(n3561), .C(n3373), .Y(n3378) );
  AOI22X1 U4176 ( .A(inst_register_registers[146]), .B(n3031), .C(
        inst_register_registers[50]), .D(n3032), .Y(n3376) );
  AOI22X1 U4177 ( .A(inst_register_registers[210]), .B(n3038), .C(
        inst_register_registers[178]), .D(n3559), .Y(n3375) );
  AOI22X1 U4178 ( .A(inst_register_registers[114]), .B(n2808), .C(
        inst_register_registers[18]), .D(n3562), .Y(n3374) );
  NAND3X1 U4179 ( .A(n3376), .B(n3375), .C(n3374), .Y(n3377) );
  OAI21X1 U4180 ( .A(n3378), .B(n3377), .C(n2795), .Y(n3379) );
  MUX2X1 U4181 ( .B(alu_result_WB[30]), .A(mem_read_data_WB[30]), .S(n3534), 
        .Y(n5231) );
  AOI22X1 U4182 ( .A(n2803), .B(inst_register_registers[30]), .C(n2802), .D(
        inst_register_registers[158]), .Y(n3380) );
  OAI21X1 U4183 ( .A(n5231), .B(n3537), .C(n3380), .Y(n3386) );
  AOI22X1 U4184 ( .A(n3207), .B(inst_register_registers[126]), .C(n3552), .D(
        inst_register_registers[254]), .Y(n3384) );
  AOI22X1 U4185 ( .A(n2807), .B(inst_register_registers[222]), .C(n2801), .D(
        inst_register_registers[190]), .Y(n3383) );
  AOI22X1 U4186 ( .A(n2805), .B(inst_register_registers[94]), .C(n2804), .D(
        inst_register_registers[62]), .Y(n3382) );
  NAND3X1 U4187 ( .A(n3384), .B(n3383), .C(n3382), .Y(n3385) );
  OAI21X1 U4188 ( .A(n3386), .B(n3385), .C(n2795), .Y(n3387) );
  AOI22X1 U4189 ( .A(n2803), .B(inst_register_registers[15]), .C(n3156), .D(
        inst_register_registers[239]), .Y(n3388) );
  OAI21X1 U4190 ( .A(n3389), .B(n3537), .C(n3388), .Y(n3394) );
  AOI22X1 U4191 ( .A(n2802), .B(inst_register_registers[143]), .C(n2804), .D(
        inst_register_registers[47]), .Y(n3392) );
  AOI22X1 U4192 ( .A(n2805), .B(inst_register_registers[79]), .C(n3535), .D(
        inst_register_registers[111]), .Y(n3391) );
  AOI22X1 U4193 ( .A(n2807), .B(inst_register_registers[207]), .C(n2801), .D(
        inst_register_registers[175]), .Y(n3390) );
  NAND3X1 U4194 ( .A(n3392), .B(n3391), .C(n3390), .Y(n3393) );
  OAI21X1 U4195 ( .A(n3394), .B(n3393), .C(n2795), .Y(n3395) );
  AOI22X1 U4196 ( .A(n2805), .B(inst_register_registers[69]), .C(n2803), .D(
        inst_register_registers[5]), .Y(n3396) );
  OAI21X1 U4197 ( .A(n5138), .B(n3148), .C(n3396), .Y(n3401) );
  AOI22X1 U4198 ( .A(n3207), .B(inst_register_registers[101]), .C(n2801), .D(
        inst_register_registers[165]), .Y(n3399) );
  AOI22X1 U4199 ( .A(n2802), .B(inst_register_registers[133]), .C(n2804), .D(
        inst_register_registers[37]), .Y(n3398) );
  AOI22X1 U4200 ( .A(n2807), .B(inst_register_registers[197]), .C(n3156), .D(
        inst_register_registers[229]), .Y(n3397) );
  NAND3X1 U4201 ( .A(n3399), .B(n3398), .C(n3397), .Y(n3400) );
  OAI21X1 U4202 ( .A(n3401), .B(n3400), .C(n2795), .Y(n3402) );
  AOI22X1 U4203 ( .A(n2805), .B(inst_register_registers[75]), .C(n2807), .D(
        inst_register_registers[203]), .Y(n3403) );
  OAI21X1 U4204 ( .A(n5156), .B(n3148), .C(n3403), .Y(n3408) );
  AOI22X1 U4205 ( .A(n2804), .B(inst_register_registers[43]), .C(n2801), .D(
        inst_register_registers[171]), .Y(n3406) );
  AOI22X1 U4206 ( .A(n3207), .B(inst_register_registers[107]), .C(n2802), .D(
        inst_register_registers[139]), .Y(n3405) );
  AOI22X1 U4207 ( .A(n2803), .B(inst_register_registers[11]), .C(n3156), .D(
        inst_register_registers[235]), .Y(n3404) );
  NAND3X1 U4208 ( .A(n3406), .B(n3405), .C(n3404), .Y(n3407) );
  OAI21X1 U4209 ( .A(n3408), .B(n3407), .C(n2795), .Y(n3409) );
  AOI22X1 U4210 ( .A(n2803), .B(inst_register_registers[8]), .C(n2801), .D(
        inst_register_registers[168]), .Y(n3410) );
  OAI21X1 U4211 ( .A(n3411), .B(n3537), .C(n3410), .Y(n3416) );
  AOI22X1 U4212 ( .A(n2805), .B(inst_register_registers[72]), .C(n2807), .D(
        inst_register_registers[200]), .Y(n3414) );
  AOI22X1 U4213 ( .A(n3207), .B(inst_register_registers[104]), .C(n2802), .D(
        inst_register_registers[136]), .Y(n3413) );
  AOI22X1 U4214 ( .A(n2804), .B(inst_register_registers[40]), .C(n3156), .D(
        inst_register_registers[232]), .Y(n3412) );
  NAND3X1 U4215 ( .A(n3414), .B(n3413), .C(n3412), .Y(n3415) );
  OAI21X1 U4216 ( .A(n3416), .B(n3415), .C(n2795), .Y(n3417) );
  AOI22X1 U4217 ( .A(inst_register_registers[252]), .B(n3073), .C(
        inst_register_registers[156]), .D(n3031), .Y(n3418) );
  OAI21X1 U4218 ( .A(n5198), .B(n3561), .C(n3418), .Y(n3424) );
  AOI22X1 U4219 ( .A(inst_register_registers[92]), .B(n2806), .C(
        inst_register_registers[220]), .D(n3419), .Y(n3422) );
  AOI22X1 U4220 ( .A(inst_register_registers[124]), .B(n2808), .C(
        inst_register_registers[60]), .D(n3563), .Y(n3421) );
  AOI22X1 U4221 ( .A(inst_register_registers[28]), .B(n3041), .C(
        inst_register_registers[188]), .D(n3559), .Y(n3420) );
  NAND3X1 U4222 ( .A(n3422), .B(n3421), .C(n3420), .Y(n3423) );
  OAI21X1 U4223 ( .A(n3424), .B(n3423), .C(n2795), .Y(n3425) );
  AOI22X1 U4224 ( .A(n2805), .B(inst_register_registers[71]), .C(n3156), .D(
        inst_register_registers[231]), .Y(n3426) );
  OAI21X1 U4225 ( .A(n5144), .B(n3148), .C(n3426), .Y(n3431) );
  AOI22X1 U4226 ( .A(n3207), .B(inst_register_registers[103]), .C(n2802), .D(
        inst_register_registers[135]), .Y(n3429) );
  AOI22X1 U4227 ( .A(n2807), .B(inst_register_registers[199]), .C(n2801), .D(
        inst_register_registers[167]), .Y(n3428) );
  AOI22X1 U4228 ( .A(n2803), .B(inst_register_registers[7]), .C(n2804), .D(
        inst_register_registers[39]), .Y(n3427) );
  NAND3X1 U4229 ( .A(n3429), .B(n3428), .C(n3427), .Y(n3430) );
  OAI21X1 U4230 ( .A(n3431), .B(n3430), .C(n2795), .Y(n3432) );
  AOI22X1 U4231 ( .A(inst_register_registers[160]), .B(n2801), .C(
        inst_register_registers[224]), .D(n3156), .Y(n3433) );
  OAI21X1 U4232 ( .A(n3434), .B(n3148), .C(n3433), .Y(n3439) );
  AOI22X1 U4233 ( .A(inst_register_registers[64]), .B(n2805), .C(
        inst_register_registers[0]), .D(n2803), .Y(n3437) );
  AOI22X1 U4234 ( .A(inst_register_registers[96]), .B(n3535), .C(
        inst_register_registers[192]), .D(n2807), .Y(n3436) );
  AOI22X1 U4235 ( .A(inst_register_registers[128]), .B(n2802), .C(
        inst_register_registers[32]), .D(n2804), .Y(n3435) );
  NAND3X1 U4236 ( .A(n3437), .B(n3436), .C(n3435), .Y(n3438) );
  OAI21X1 U4237 ( .A(n3439), .B(n3438), .C(n2795), .Y(n3440) );
  AOI22X1 U4238 ( .A(n2807), .B(inst_register_registers[206]), .C(n3552), .D(
        inst_register_registers[238]), .Y(n3441) );
  OAI21X1 U4239 ( .A(n3442), .B(n3537), .C(n3441), .Y(n3447) );
  AOI22X1 U4240 ( .A(n2805), .B(inst_register_registers[78]), .C(n2802), .D(
        inst_register_registers[142]), .Y(n3445) );
  AOI22X1 U4241 ( .A(n2803), .B(inst_register_registers[14]), .C(n2801), .D(
        inst_register_registers[174]), .Y(n3444) );
  AOI22X1 U4242 ( .A(n3207), .B(inst_register_registers[110]), .C(n2804), .D(
        inst_register_registers[46]), .Y(n3443) );
  NAND3X1 U4243 ( .A(n3445), .B(n3444), .C(n3443), .Y(n3446) );
  OAI21X1 U4244 ( .A(n3447), .B(n3446), .C(n2795), .Y(n3448) );
  AOI22X1 U4245 ( .A(n2803), .B(inst_register_registers[2]), .C(n3207), .D(
        inst_register_registers[98]), .Y(n3449) );
  OAI21X1 U4246 ( .A(n5129), .B(n3148), .C(n3449), .Y(n3454) );
  AOI22X1 U4247 ( .A(n2807), .B(inst_register_registers[194]), .C(n2804), .D(
        inst_register_registers[34]), .Y(n3452) );
  AOI22X1 U4248 ( .A(n2805), .B(inst_register_registers[66]), .C(n3156), .D(
        inst_register_registers[226]), .Y(n3451) );
  AOI22X1 U4249 ( .A(n2802), .B(inst_register_registers[130]), .C(n2801), .D(
        inst_register_registers[162]), .Y(n3450) );
  NAND3X1 U4250 ( .A(n3452), .B(n3451), .C(n3450), .Y(n3453) );
  OAI21X1 U4251 ( .A(n3454), .B(n3453), .C(n2795), .Y(n3455) );
  AOI22X1 U4252 ( .A(n2805), .B(inst_register_registers[83]), .C(n2802), .D(
        inst_register_registers[147]), .Y(n3456) );
  OAI21X1 U4253 ( .A(n3652), .B(n3148), .C(n3456), .Y(n3461) );
  AOI22X1 U4254 ( .A(n2803), .B(inst_register_registers[19]), .C(n2804), .D(
        inst_register_registers[51]), .Y(n3459) );
  AOI22X1 U4255 ( .A(n2801), .B(inst_register_registers[179]), .C(n3552), .D(
        inst_register_registers[243]), .Y(n3458) );
  AOI22X1 U4256 ( .A(n3207), .B(inst_register_registers[115]), .C(n2807), .D(
        inst_register_registers[211]), .Y(n3457) );
  NAND3X1 U4257 ( .A(n3459), .B(n3458), .C(n3457), .Y(n3460) );
  OAI21X1 U4258 ( .A(n3461), .B(n3460), .C(n2795), .Y(n3462) );
  AOI22X1 U4259 ( .A(n2805), .B(inst_register_registers[74]), .C(n2803), .D(
        inst_register_registers[10]), .Y(n3463) );
  OAI21X1 U4260 ( .A(n5152), .B(n3537), .C(n3463), .Y(n3468) );
  AOI22X1 U4261 ( .A(n2804), .B(inst_register_registers[42]), .C(n3156), .D(
        inst_register_registers[234]), .Y(n3466) );
  AOI22X1 U4262 ( .A(n2802), .B(inst_register_registers[138]), .C(n2801), .D(
        inst_register_registers[170]), .Y(n3465) );
  AOI22X1 U4263 ( .A(n3207), .B(inst_register_registers[106]), .C(n2807), .D(
        inst_register_registers[202]), .Y(n3464) );
  NAND3X1 U4264 ( .A(n3466), .B(n3465), .C(n3464), .Y(n3467) );
  OAI21X1 U4265 ( .A(n3468), .B(n3467), .C(n2795), .Y(n3469) );
  AOI22X1 U4266 ( .A(n2803), .B(inst_register_registers[12]), .C(n3156), .D(
        inst_register_registers[236]), .Y(n3470) );
  OAI21X1 U4267 ( .A(n5159), .B(n3148), .C(n3470), .Y(n3475) );
  AOI22X1 U4268 ( .A(n3207), .B(inst_register_registers[108]), .C(n2802), .D(
        inst_register_registers[140]), .Y(n3473) );
  AOI22X1 U4269 ( .A(n2804), .B(inst_register_registers[44]), .C(n2801), .D(
        inst_register_registers[172]), .Y(n3472) );
  AOI22X1 U4270 ( .A(n2805), .B(inst_register_registers[76]), .C(n2807), .D(
        inst_register_registers[204]), .Y(n3471) );
  NAND3X1 U4271 ( .A(n3473), .B(n3472), .C(n3471), .Y(n3474) );
  OAI21X1 U4272 ( .A(n3475), .B(n3474), .C(n2795), .Y(n3476) );
  AOI22X1 U4273 ( .A(n3207), .B(inst_register_registers[102]), .C(n2804), .D(
        inst_register_registers[38]), .Y(n3477) );
  OAI21X1 U4274 ( .A(n5141), .B(n3148), .C(n3477), .Y(n3482) );
  AOI22X1 U4275 ( .A(n2803), .B(inst_register_registers[6]), .C(n2801), .D(
        inst_register_registers[166]), .Y(n3480) );
  AOI22X1 U4276 ( .A(n2805), .B(inst_register_registers[70]), .C(n2802), .D(
        inst_register_registers[134]), .Y(n3479) );
  AOI22X1 U4277 ( .A(n2807), .B(inst_register_registers[198]), .C(n3156), .D(
        inst_register_registers[230]), .Y(n3478) );
  NAND3X1 U4278 ( .A(n3480), .B(n3479), .C(n3478), .Y(n3481) );
  OAI21X1 U4279 ( .A(n3482), .B(n3481), .C(n2795), .Y(n3483) );
  AOI22X1 U4280 ( .A(n2802), .B(inst_register_registers[131]), .C(n2804), .D(
        inst_register_registers[35]), .Y(n3484) );
  OAI21X1 U4281 ( .A(n5132), .B(n3148), .C(n3484), .Y(n3489) );
  AOI22X1 U4282 ( .A(n2801), .B(inst_register_registers[163]), .C(n3156), .D(
        inst_register_registers[227]), .Y(n3487) );
  AOI22X1 U4283 ( .A(n2805), .B(inst_register_registers[67]), .C(n2803), .D(
        inst_register_registers[3]), .Y(n3486) );
  AOI22X1 U4284 ( .A(n3207), .B(inst_register_registers[99]), .C(n2807), .D(
        inst_register_registers[195]), .Y(n3485) );
  NAND3X1 U4285 ( .A(n3487), .B(n3486), .C(n3485), .Y(n3488) );
  OAI21X1 U4286 ( .A(n3489), .B(n3488), .C(n2795), .Y(n3490) );
  AOI22X1 U4287 ( .A(n2807), .B(inst_register_registers[209]), .C(n2804), .D(
        inst_register_registers[49]), .Y(n3491) );
  OAI21X1 U4288 ( .A(n5171), .B(n3148), .C(n3491), .Y(n3496) );
  AOI22X1 U4289 ( .A(n2803), .B(inst_register_registers[17]), .C(n3535), .D(
        inst_register_registers[113]), .Y(n3494) );
  AOI22X1 U4290 ( .A(n2805), .B(inst_register_registers[81]), .C(n3552), .D(
        inst_register_registers[241]), .Y(n3493) );
  AOI22X1 U4291 ( .A(n2802), .B(inst_register_registers[145]), .C(n2801), .D(
        inst_register_registers[177]), .Y(n3492) );
  NAND3X1 U4292 ( .A(n3494), .B(n3493), .C(n3492), .Y(n3495) );
  OAI21X1 U4293 ( .A(n3496), .B(n3495), .C(n2795), .Y(n3497) );
  AOI22X1 U4294 ( .A(n2804), .B(inst_register_registers[50]), .C(n2801), .D(
        inst_register_registers[178]), .Y(n3498) );
  OAI21X1 U4295 ( .A(n3656), .B(n3537), .C(n3498), .Y(n3503) );
  AOI22X1 U4296 ( .A(n3207), .B(inst_register_registers[114]), .C(n2807), .D(
        inst_register_registers[210]), .Y(n3501) );
  AOI22X1 U4297 ( .A(n2803), .B(inst_register_registers[18]), .C(n2802), .D(
        inst_register_registers[146]), .Y(n3500) );
  AOI22X1 U4298 ( .A(n2805), .B(inst_register_registers[82]), .C(n3156), .D(
        inst_register_registers[242]), .Y(n3499) );
  NAND3X1 U4299 ( .A(n3501), .B(n3500), .C(n3499), .Y(n3502) );
  OAI21X1 U4300 ( .A(n3503), .B(n3502), .C(n2795), .Y(n3504) );
  AOI22X1 U4301 ( .A(n2805), .B(inst_register_registers[80]), .C(n2803), .D(
        inst_register_registers[16]), .Y(n3505) );
  OAI21X1 U4302 ( .A(n3506), .B(n3537), .C(n3505), .Y(n3511) );
  AOI22X1 U4303 ( .A(n3207), .B(inst_register_registers[112]), .C(n3552), .D(
        inst_register_registers[240]), .Y(n3509) );
  AOI22X1 U4304 ( .A(n2802), .B(inst_register_registers[144]), .C(n2801), .D(
        inst_register_registers[176]), .Y(n3508) );
  AOI22X1 U4305 ( .A(n2807), .B(inst_register_registers[208]), .C(n2804), .D(
        inst_register_registers[48]), .Y(n3507) );
  NAND3X1 U4306 ( .A(n3509), .B(n3508), .C(n3507), .Y(n3510) );
  OAI21X1 U4307 ( .A(n3511), .B(n3510), .C(n2795), .Y(n3512) );
  AOI22X1 U4308 ( .A(n2803), .B(inst_register_registers[1]), .C(n2807), .D(
        inst_register_registers[193]), .Y(n3513) );
  OAI21X1 U4309 ( .A(n5126), .B(n3148), .C(n3513), .Y(n3518) );
  AOI22X1 U4310 ( .A(n2801), .B(inst_register_registers[161]), .C(n3156), .D(
        inst_register_registers[225]), .Y(n3516) );
  AOI22X1 U4311 ( .A(n2805), .B(inst_register_registers[65]), .C(n2802), .D(
        inst_register_registers[129]), .Y(n3515) );
  AOI22X1 U4312 ( .A(n3207), .B(inst_register_registers[97]), .C(n2804), .D(
        inst_register_registers[33]), .Y(n3514) );
  NAND3X1 U4313 ( .A(n3516), .B(n3515), .C(n3514), .Y(n3517) );
  OAI21X1 U4314 ( .A(n3518), .B(n3517), .C(n2795), .Y(n3519) );
  AOI22X1 U4315 ( .A(n2803), .B(inst_register_registers[9]), .C(n2802), .D(
        inst_register_registers[137]), .Y(n3520) );
  OAI21X1 U4316 ( .A(n5149), .B(n3537), .C(n3520), .Y(n3525) );
  AOI22X1 U4317 ( .A(n2805), .B(inst_register_registers[73]), .C(n3535), .D(
        inst_register_registers[105]), .Y(n3523) );
  AOI22X1 U4318 ( .A(n2801), .B(inst_register_registers[169]), .C(n3156), .D(
        inst_register_registers[233]), .Y(n3522) );
  AOI22X1 U4319 ( .A(n2807), .B(inst_register_registers[201]), .C(n2804), .D(
        inst_register_registers[41]), .Y(n3521) );
  NAND3X1 U4320 ( .A(n3523), .B(n3522), .C(n3521), .Y(n3524) );
  OAI21X1 U4321 ( .A(n3525), .B(n3524), .C(n2795), .Y(n3526) );
  AOI22X1 U4322 ( .A(n2803), .B(inst_register_registers[4]), .C(n2807), .D(
        inst_register_registers[196]), .Y(n3527) );
  OAI21X1 U4323 ( .A(n5135), .B(n3148), .C(n3527), .Y(n3532) );
  AOI22X1 U4324 ( .A(n2804), .B(inst_register_registers[36]), .C(n2801), .D(
        inst_register_registers[164]), .Y(n3530) );
  AOI22X1 U4325 ( .A(n3207), .B(inst_register_registers[100]), .C(n3156), .D(
        inst_register_registers[228]), .Y(n3529) );
  AOI22X1 U4326 ( .A(n2805), .B(inst_register_registers[68]), .C(n2802), .D(
        inst_register_registers[132]), .Y(n3528) );
  NAND3X1 U4327 ( .A(n3530), .B(n3529), .C(n3528), .Y(n3531) );
  OAI21X1 U4328 ( .A(n3532), .B(n3531), .C(n2795), .Y(n3533) );
  MUX2X1 U4329 ( .B(alu_result_WB[29]), .A(mem_read_data_WB[29]), .S(n3534), 
        .Y(n5121) );
  AOI22X1 U4330 ( .A(n3535), .B(inst_register_registers[125]), .C(n3552), .D(
        inst_register_registers[253]), .Y(n3536) );
  OAI21X1 U4331 ( .A(n5121), .B(n3537), .C(n3536), .Y(n3542) );
  AOI22X1 U4332 ( .A(n2803), .B(inst_register_registers[29]), .C(n2801), .D(
        inst_register_registers[189]), .Y(n3540) );
  AOI22X1 U4333 ( .A(n2805), .B(inst_register_registers[93]), .C(n2802), .D(
        inst_register_registers[157]), .Y(n3539) );
  AOI22X1 U4334 ( .A(n2807), .B(inst_register_registers[221]), .C(n2804), .D(
        inst_register_registers[61]), .Y(n3538) );
  NAND3X1 U4335 ( .A(n3540), .B(n3539), .C(n3538), .Y(n3541) );
  OAI21X1 U4336 ( .A(n3542), .B(n3541), .C(n2795), .Y(n3543) );
  AOI22X1 U4337 ( .A(inst_register_registers[253]), .B(n3073), .C(
        inst_register_registers[125]), .D(n2808), .Y(n3544) );
  OAI21X1 U4338 ( .A(n5121), .B(n3561), .C(n3544), .Y(n3549) );
  AOI22X1 U4339 ( .A(inst_register_registers[29]), .B(n3041), .C(
        inst_register_registers[221]), .D(n3038), .Y(n3547) );
  AOI22X1 U4340 ( .A(inst_register_registers[189]), .B(n3071), .C(
        inst_register_registers[157]), .D(n3564), .Y(n3546) );
  AOI22X1 U4341 ( .A(inst_register_registers[93]), .B(n2806), .C(
        inst_register_registers[61]), .D(n3563), .Y(n3545) );
  NAND3X1 U4342 ( .A(n3547), .B(n3546), .C(n3545), .Y(n3548) );
  OAI21X1 U4343 ( .A(n3549), .B(n3548), .C(n2795), .Y(n3550) );
  AOI22X1 U4344 ( .A(n2803), .B(inst_register_registers[13]), .C(n2804), .D(
        inst_register_registers[45]), .Y(n3551) );
  OAI21X1 U4345 ( .A(n5162), .B(n3148), .C(n3551), .Y(n3557) );
  AOI22X1 U4346 ( .A(n3207), .B(inst_register_registers[109]), .C(n3552), .D(
        inst_register_registers[237]), .Y(n3555) );
  AOI22X1 U4347 ( .A(n2807), .B(inst_register_registers[205]), .C(n2801), .D(
        inst_register_registers[173]), .Y(n3554) );
  AOI22X1 U4348 ( .A(n2805), .B(inst_register_registers[77]), .C(n2802), .D(
        inst_register_registers[141]), .Y(n3553) );
  NAND3X1 U4349 ( .A(n3555), .B(n3554), .C(n3553), .Y(n3556) );
  OAI21X1 U4350 ( .A(n3557), .B(n3556), .C(n2795), .Y(n3558) );
  AOI22X1 U4351 ( .A(inst_register_registers[190]), .B(n3559), .C(
        inst_register_registers[94]), .D(n2806), .Y(n3560) );
  OAI21X1 U4352 ( .A(n5231), .B(n3561), .C(n3560), .Y(n3569) );
  AOI22X1 U4353 ( .A(inst_register_registers[222]), .B(n3038), .C(
        inst_register_registers[30]), .D(n3562), .Y(n3567) );
  AOI22X1 U4354 ( .A(inst_register_registers[126]), .B(n2808), .C(
        inst_register_registers[62]), .D(n3563), .Y(n3566) );
  AOI22X1 U4355 ( .A(inst_register_registers[254]), .B(n3073), .C(
        inst_register_registers[158]), .D(n3564), .Y(n3565) );
  NAND3X1 U4356 ( .A(n3567), .B(n3566), .C(n3565), .Y(n3568) );
  OAI21X1 U4357 ( .A(n3569), .B(n3568), .C(n2795), .Y(n3570) );
  FAX1 U4358 ( .A(n4086), .B(n3572), .C(n3571), .YC(n3578), .YS(n3576) );
  NAND2X1 U4359 ( .A(n4086), .B(n4092), .Y(n3574) );
  OAI21X1 U4360 ( .A(n4092), .B(n4086), .C(n3739), .Y(n3573) );
  OAI21X1 U4361 ( .A(n3574), .B(n3953), .C(n3573), .Y(n3575) );
  AOI21X1 U4362 ( .A(n4263), .B(n3576), .C(n3575), .Y(n3577) );
  FAX1 U4363 ( .A(n4089), .B(n3579), .C(n3578), .YC(n3585), .YS(n3583) );
  NAND2X1 U4364 ( .A(n4089), .B(n4090), .Y(n3581) );
  OAI21X1 U4365 ( .A(n4090), .B(n4089), .C(n3739), .Y(n3580) );
  OAI21X1 U4366 ( .A(n3581), .B(n3953), .C(n3580), .Y(n3582) );
  AOI21X1 U4367 ( .A(n4263), .B(n3583), .C(n3582), .Y(n3584) );
  FAX1 U4368 ( .A(n4095), .B(n3586), .C(n3585), .YC(n3007), .YS(n3590) );
  NAND2X1 U4369 ( .A(n4095), .B(n4098), .Y(n3588) );
  OAI21X1 U4370 ( .A(n4098), .B(n4095), .C(n3739), .Y(n3587) );
  OAI21X1 U4371 ( .A(n3588), .B(n4047), .C(n3587), .Y(n3589) );
  AOI21X1 U4372 ( .A(n4263), .B(n3590), .C(n3589), .Y(n3591) );
  NOR2X1 U4373 ( .A(n4434), .B(n4432), .Y(n4439) );
  NAND2X1 U4374 ( .A(alu_result_MEM[0]), .B(n4439), .Y(n4433) );
  INVX1 U4375 ( .A(n3592), .Y(n3593) );
  INVX1 U4376 ( .A(op_type_MEM[3]), .Y(n3767) );
  NAND2X1 U4377 ( .A(n3593), .B(n3767), .Y(n3594) );
  OAI21X1 U4378 ( .A(n4433), .B(n3594), .C(n2815), .Y(n5061) );
  INVX2 U4379 ( .A(n5009), .Y(n5065) );
  INVX1 U4380 ( .A(n4433), .Y(n3595) );
  NAND2X1 U4381 ( .A(n3595), .B(n4927), .Y(n3596) );
  OAI22X1 U4382 ( .A(inst_data_MEM_data[227]), .B(n5065), .C(
        write_mem_data_MEM[3]), .D(n5014), .Y(n3597) );
  AND2X2 U4383 ( .A(n4426), .B(shifted_address_EX[0]), .Y(inst_EX2MEM_reg_N7)
         );
  AND2X2 U4384 ( .A(n4426), .B(shifted_address_EX[1]), .Y(inst_EX2MEM_reg_N8)
         );
  NOR2X1 U4385 ( .A(jump_inst_addr_EX[0]), .B(inst_addr_EX[2]), .Y(n3598) );
  NAND2X1 U4386 ( .A(n3598), .B(n3766), .Y(n4333) );
  NOR2X1 U4387 ( .A(n3598), .B(n3766), .Y(n4335) );
  AOI21X1 U4388 ( .A(inst_addr_EX[3]), .B(n4333), .C(n4335), .Y(n3599) );
  NAND2X1 U4389 ( .A(n3599), .B(n3765), .Y(n4338) );
  NOR2X1 U4390 ( .A(n3599), .B(n3765), .Y(n4340) );
  AOI21X1 U4391 ( .A(inst_addr_EX[4]), .B(n4338), .C(n4340), .Y(n3600) );
  NAND2X1 U4392 ( .A(n3600), .B(n3764), .Y(n4343) );
  NOR2X1 U4393 ( .A(n3600), .B(n3764), .Y(n4345) );
  AOI21X1 U4394 ( .A(inst_addr_EX[5]), .B(n4343), .C(n4345), .Y(n3601) );
  NAND2X1 U4395 ( .A(n3601), .B(n3763), .Y(n4348) );
  NOR2X1 U4396 ( .A(n3601), .B(n3763), .Y(n4350) );
  AOI21X1 U4397 ( .A(inst_addr_EX[6]), .B(n4348), .C(n4350), .Y(n3602) );
  NAND2X1 U4398 ( .A(n3602), .B(n3762), .Y(n4353) );
  NOR2X1 U4399 ( .A(n3602), .B(n3762), .Y(n4355) );
  AOI21X1 U4400 ( .A(inst_addr_EX[7]), .B(n4353), .C(n4355), .Y(n3604) );
  INVX1 U4401 ( .A(n3604), .Y(n3603) );
  NOR2X1 U4402 ( .A(jump_inst_addr_EX[6]), .B(n3603), .Y(n4358) );
  INVX1 U4403 ( .A(inst_addr_EX[8]), .Y(n3606) );
  NOR2X1 U4404 ( .A(n3604), .B(n3761), .Y(n4359) );
  INVX1 U4405 ( .A(n4359), .Y(n3605) );
  OAI21X1 U4406 ( .A(n4358), .B(n3606), .C(n3605), .Y(n3608) );
  AND2X2 U4407 ( .A(n4426), .B(n3607), .Y(inst_EX2MEM_reg_N16) );
  FAX1 U4408 ( .A(inst_addr_EX[9]), .B(jump_inst_addr_EX[7]), .C(n3608), .YC(
        n4363), .YS(n3607) );
  NOR2X1 U4409 ( .A(jump_inst_addr_EX[8]), .B(n4363), .Y(n4362) );
  INVX1 U4410 ( .A(inst_addr_EX[10]), .Y(n3610) );
  NAND2X1 U4411 ( .A(jump_inst_addr_EX[8]), .B(n4363), .Y(n3609) );
  OAI21X1 U4412 ( .A(n4362), .B(n3610), .C(n3609), .Y(n4366) );
  INVX1 U4413 ( .A(n4366), .Y(n3612) );
  OAI21X1 U4414 ( .A(jump_inst_addr_EX[9]), .B(n4366), .C(inst_addr_EX[11]), 
        .Y(n3611) );
  OAI21X1 U4415 ( .A(n3612), .B(n4367), .C(n3611), .Y(n3614) );
  AND2X2 U4416 ( .A(n4426), .B(n3613), .Y(inst_EX2MEM_reg_N19) );
  FAX1 U4417 ( .A(inst_addr_EX[12]), .B(jump_inst_addr_EX[10]), .C(n3614), 
        .YC(n4371), .YS(n3613) );
  NOR2X1 U4418 ( .A(jump_inst_addr_EX[11]), .B(n4371), .Y(n4370) );
  INVX1 U4419 ( .A(inst_addr_EX[13]), .Y(n3616) );
  NAND2X1 U4420 ( .A(jump_inst_addr_EX[11]), .B(n4371), .Y(n3615) );
  OAI21X1 U4421 ( .A(n4370), .B(n3616), .C(n3615), .Y(n4374) );
  INVX1 U4422 ( .A(n4374), .Y(n3618) );
  OAI21X1 U4423 ( .A(jump_inst_addr_EX[12]), .B(n4374), .C(inst_addr_EX[14]), 
        .Y(n3617) );
  OAI21X1 U4424 ( .A(n3618), .B(n4375), .C(n3617), .Y(n3620) );
  AND2X2 U4425 ( .A(n4426), .B(n3619), .Y(inst_EX2MEM_reg_N22) );
  FAX1 U4426 ( .A(inst_addr_EX[15]), .B(jump_inst_addr_EX[13]), .C(n3620), 
        .YC(n4379), .YS(n3619) );
  NOR2X1 U4427 ( .A(jump_inst_addr_EX[14]), .B(n4379), .Y(n4378) );
  INVX1 U4428 ( .A(inst_addr_EX[16]), .Y(n3622) );
  NAND2X1 U4429 ( .A(jump_inst_addr_EX[14]), .B(n4379), .Y(n3621) );
  OAI21X1 U4430 ( .A(n4378), .B(n3622), .C(n3621), .Y(n4382) );
  INVX1 U4431 ( .A(n4382), .Y(n3624) );
  OAI21X1 U4432 ( .A(n4414), .B(n4382), .C(inst_addr_EX[17]), .Y(n3623) );
  OAI21X1 U4433 ( .A(n3624), .B(n4419), .C(n3623), .Y(n3626) );
  AND2X2 U4434 ( .A(n4426), .B(n3625), .Y(inst_EX2MEM_reg_N25) );
  FAX1 U4435 ( .A(inst_addr_EX[18]), .B(n4414), .C(n3626), .YC(n4386), .YS(
        n3625) );
  NOR2X1 U4436 ( .A(n4414), .B(n4386), .Y(n4385) );
  NAND2X1 U4437 ( .A(n4414), .B(n4386), .Y(n3627) );
  OAI21X1 U4438 ( .A(n4385), .B(n3628), .C(n3627), .Y(n3640) );
  AND2X2 U4439 ( .A(n4426), .B(n3629), .Y(inst_EX2MEM_reg_N27) );
  NAND2X1 U4440 ( .A(inst_address[13]), .B(inst_address[12]), .Y(n3846) );
  INVX1 U4441 ( .A(inst_address[3]), .Y(n4742) );
  INVX1 U4442 ( .A(inst_address[2]), .Y(n5502) );
  NOR2X1 U4443 ( .A(n4742), .B(n5502), .Y(n3934) );
  NAND2X1 U4444 ( .A(n3934), .B(inst_address[4]), .Y(n4273) );
  INVX1 U4445 ( .A(inst_address[5]), .Y(n4738) );
  NOR2X1 U4446 ( .A(n4273), .B(n4738), .Y(n4280) );
  NAND2X1 U4447 ( .A(n4280), .B(inst_address[6]), .Y(n4279) );
  INVX1 U4448 ( .A(inst_address[7]), .Y(n4734) );
  NOR2X1 U4449 ( .A(n4279), .B(n4734), .Y(n3924) );
  NAND3X1 U4450 ( .A(n3924), .B(inst_address[9]), .C(inst_address[8]), .Y(
        n3913) );
  INVX1 U4451 ( .A(inst_address[10]), .Y(n4728) );
  NOR2X1 U4452 ( .A(n3913), .B(n4728), .Y(n3909) );
  NAND2X1 U4453 ( .A(n3909), .B(inst_address[11]), .Y(n3854) );
  NAND2X1 U4454 ( .A(n2795), .B(n3632), .Y(n4286) );
  NAND2X1 U4455 ( .A(n3633), .B(n4290), .Y(n3630) );
  NOR2X1 U4456 ( .A(inst_address[14]), .B(n3630), .Y(n3851) );
  INVX2 U4457 ( .A(n2795), .Y(n5524) );
  NOR2X1 U4458 ( .A(n5392), .B(n3631), .Y(n4617) );
  NOR2X1 U4459 ( .A(n3632), .B(n3933), .Y(n3908) );
  NOR2X1 U4460 ( .A(n4617), .B(n3908), .Y(n4289) );
  OAI21X1 U4461 ( .A(n3633), .B(n5524), .C(n4289), .Y(n3850) );
  INVX1 U4462 ( .A(inst_address[14]), .Y(n4719) );
  INVX1 U4463 ( .A(n3634), .Y(n3635) );
  NOR2X1 U4464 ( .A(n3635), .B(n2796), .Y(n5526) );
  INVX2 U4465 ( .A(n4305), .Y(n4294) );
  NOR2X1 U4466 ( .A(n3637), .B(n2796), .Y(n3902) );
  BUFX2 U4467 ( .A(n3902), .Y(n5497) );
  AOI22X1 U4468 ( .A(n4294), .B(shifted_address_MEM[14]), .C(n5497), .D(
        jump_inst_addr_MEM[14]), .Y(n3638) );
  OAI21X1 U4469 ( .A(n4293), .B(n4719), .C(n3638), .Y(n3639) );
  FAX1 U4470 ( .A(inst_addr_EX[20]), .B(n4414), .C(n3640), .YC(n4390), .YS(
        n3629) );
  AOI21X1 U4471 ( .A(inst_addr_EX[21]), .B(n4390), .C(n4414), .Y(n4394) );
  INVX1 U4472 ( .A(inst_addr_EX[22]), .Y(n3641) );
  OAI21X1 U4473 ( .A(n4394), .B(n3641), .C(n4419), .Y(n4399) );
  INVX1 U4474 ( .A(inst_addr_EX[23]), .Y(n3642) );
  INVX1 U4475 ( .A(inst_addr_EX[21]), .Y(n4393) );
  NAND2X1 U4476 ( .A(n4414), .B(n4390), .Y(n4389) );
  NAND2X1 U4477 ( .A(n4393), .B(n4389), .Y(n4395) );
  OAI21X1 U4478 ( .A(inst_addr_EX[22]), .B(n4395), .C(n4414), .Y(n4398) );
  OAI21X1 U4479 ( .A(n3643), .B(n3642), .C(n4398), .Y(n3645) );
  AND2X2 U4480 ( .A(n4426), .B(n3644), .Y(inst_EX2MEM_reg_N31) );
  FAX1 U4481 ( .A(inst_addr_EX[24]), .B(n4414), .C(n3645), .YC(n3647), .YS(
        n3644) );
  AND2X2 U4482 ( .A(n4426), .B(n3646), .Y(inst_EX2MEM_reg_N32) );
  FAX1 U4483 ( .A(inst_addr_EX[25]), .B(n4414), .C(n3647), .YC(n4403), .YS(
        n3646) );
  AOI21X1 U4484 ( .A(inst_addr_EX[26]), .B(n4403), .C(n4414), .Y(n4408) );
  INVX1 U4485 ( .A(inst_addr_EX[27]), .Y(n3649) );
  INVX1 U4486 ( .A(inst_addr_EX[26]), .Y(n4406) );
  NAND2X1 U4487 ( .A(n4414), .B(n4403), .Y(n4402) );
  AOI21X1 U4488 ( .A(n4406), .B(n4402), .C(n4419), .Y(n4407) );
  INVX1 U4489 ( .A(n4407), .Y(n3648) );
  OAI21X1 U4490 ( .A(n4408), .B(n3649), .C(n3648), .Y(n4411) );
  AND2X2 U4491 ( .A(n4426), .B(n3650), .Y(inst_EX2MEM_reg_N35) );
  AOI22X1 U4492 ( .A(reg_read_data_1_EX[19]), .B(n3947), .C(alu_result_MEM[19]), .D(n2814), .Y(n3651) );
  OAI21X1 U4493 ( .A(n3652), .B(n3733), .C(n3651), .Y(n4062) );
  AOI22X1 U4494 ( .A(n3941), .B(reg_read_data_2_EX[19]), .C(alu_result_MEM[19]), .D(n3942), .Y(n3654) );
  NAND2X1 U4495 ( .A(n5176), .B(n3946), .Y(n3653) );
  NAND3X1 U4496 ( .A(n3943), .B(n3654), .C(n3653), .Y(n4058) );
  XOR2X1 U4497 ( .A(n4259), .B(n4058), .Y(n3678) );
  AOI22X1 U4498 ( .A(reg_read_data_1_EX[18]), .B(n3947), .C(alu_result_MEM[18]), .D(n2814), .Y(n3655) );
  OAI21X1 U4499 ( .A(n3656), .B(n3733), .C(n3655), .Y(n4138) );
  AOI22X1 U4500 ( .A(alu_result_MEM[18]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[18]), .Y(n3657) );
  NAND2X1 U4501 ( .A(n3657), .B(n3943), .Y(n3658) );
  AOI21X1 U4502 ( .A(n5174), .B(n3946), .C(n3658), .Y(n4139) );
  XOR2X1 U4503 ( .A(n4259), .B(n4056), .Y(n4005) );
  AOI22X1 U4504 ( .A(reg_read_data_1_EX[17]), .B(n3947), .C(alu_result_MEM[17]), .D(n2814), .Y(n3659) );
  OAI21X1 U4505 ( .A(n5171), .B(n3733), .C(n3659), .Y(n4063) );
  AOI22X1 U4506 ( .A(alu_result_MEM[17]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[17]), .Y(n3660) );
  AND2X2 U4507 ( .A(n3943), .B(n3660), .Y(n3661) );
  OAI21X1 U4508 ( .A(n5171), .B(n3736), .C(n3661), .Y(n4135) );
  XOR2X1 U4509 ( .A(n4259), .B(n4135), .Y(n4012) );
  FAX1 U4510 ( .A(n4112), .B(n3663), .C(n3662), .YC(n4011), .YS(n2977) );
  NAND2X1 U4511 ( .A(n4062), .B(n4058), .Y(n3665) );
  OAI21X1 U4512 ( .A(n4062), .B(n4058), .C(n3739), .Y(n3664) );
  OAI21X1 U4513 ( .A(n3665), .B(n4047), .C(n3664), .Y(n3666) );
  AOI21X1 U4514 ( .A(n4263), .B(n3667), .C(n3666), .Y(n3668) );
  INVX1 U4515 ( .A(n3668), .Y(inst_EX2MEM_reg_N58) );
  AOI22X1 U4516 ( .A(reg_read_data_1_EX[21]), .B(n3947), .C(alu_result_MEM[21]), .D(n2814), .Y(n3669) );
  OAI21X1 U4517 ( .A(n3670), .B(n3733), .C(n3669), .Y(n4144) );
  AOI22X1 U4518 ( .A(alu_result_MEM[21]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[21]), .Y(n3672) );
  NAND2X1 U4519 ( .A(n5180), .B(n3946), .Y(n3671) );
  NAND3X1 U4520 ( .A(n3943), .B(n3672), .C(n3671), .Y(n4054) );
  XOR2X1 U4521 ( .A(n4259), .B(n4054), .Y(n3689) );
  AOI22X1 U4522 ( .A(reg_read_data_1_EX[20]), .B(n3947), .C(alu_result_MEM[20]), .D(n2814), .Y(n3673) );
  OAI21X1 U4523 ( .A(n3674), .B(n3733), .C(n3673), .Y(n4060) );
  AOI22X1 U4524 ( .A(alu_result_MEM[20]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[20]), .Y(n3675) );
  NAND2X1 U4525 ( .A(n3675), .B(n3943), .Y(n3676) );
  AOI21X1 U4526 ( .A(n5178), .B(n3946), .C(n3676), .Y(n4059) );
  XOR2X1 U4527 ( .A(n4259), .B(n4001), .Y(n3997) );
  FAX1 U4528 ( .A(n4062), .B(n3678), .C(n3677), .YC(n3996), .YS(n3667) );
  NAND2X1 U4529 ( .A(n4144), .B(n4054), .Y(n3680) );
  OAI21X1 U4530 ( .A(n4144), .B(n4054), .C(n3739), .Y(n3679) );
  OAI21X1 U4531 ( .A(n3680), .B(n3953), .C(n3679), .Y(n3681) );
  AOI21X1 U4532 ( .A(n4263), .B(n3682), .C(n3681), .Y(n3683) );
  INVX1 U4533 ( .A(n3683), .Y(inst_EX2MEM_reg_N60) );
  AOI22X1 U4534 ( .A(reg_read_data_1_EX[22]), .B(n3947), .C(alu_result_MEM[22]), .D(n2814), .Y(n3684) );
  OAI21X1 U4535 ( .A(n3685), .B(n3733), .C(n3684), .Y(n4146) );
  AOI22X1 U4536 ( .A(alu_result_MEM[22]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[22]), .Y(n3687) );
  NAND2X1 U4537 ( .A(n5182), .B(n3946), .Y(n3686) );
  NAND3X1 U4538 ( .A(n3943), .B(n3687), .C(n3686), .Y(n4143) );
  XOR2X1 U4539 ( .A(n4259), .B(n4143), .Y(n3700) );
  FAX1 U4540 ( .A(n4144), .B(n3689), .C(n3688), .YC(n3699), .YS(n3682) );
  NAND2X1 U4541 ( .A(n4146), .B(n4143), .Y(n3691) );
  OAI21X1 U4542 ( .A(n4146), .B(n4143), .C(n3739), .Y(n3690) );
  OAI21X1 U4543 ( .A(n3691), .B(n3953), .C(n3690), .Y(n3692) );
  AOI21X1 U4544 ( .A(n4263), .B(n3693), .C(n3692), .Y(n3694) );
  INVX1 U4545 ( .A(n3694), .Y(inst_EX2MEM_reg_N61) );
  AOI22X1 U4546 ( .A(reg_read_data_1_EX[23]), .B(n3947), .C(alu_result_MEM[23]), .D(n2814), .Y(n3695) );
  OAI21X1 U4547 ( .A(n3696), .B(n3733), .C(n3695), .Y(n4160) );
  AOI22X1 U4548 ( .A(alu_result_MEM[23]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[23]), .Y(n3698) );
  NAND2X1 U4549 ( .A(n5184), .B(n3946), .Y(n3697) );
  NAND3X1 U4550 ( .A(n3943), .B(n3698), .C(n3697), .Y(n4157) );
  XOR2X1 U4551 ( .A(n4259), .B(n4157), .Y(n3713) );
  FAX1 U4552 ( .A(n4146), .B(n3700), .C(n3699), .YC(n3712), .YS(n3693) );
  NAND2X1 U4553 ( .A(n4160), .B(n4157), .Y(n3702) );
  OAI21X1 U4554 ( .A(n4160), .B(n4157), .C(n3739), .Y(n3701) );
  OAI21X1 U4555 ( .A(n3702), .B(n3953), .C(n3701), .Y(n3703) );
  AOI21X1 U4556 ( .A(n4263), .B(n3704), .C(n3703), .Y(n3705) );
  INVX1 U4557 ( .A(n3705), .Y(inst_EX2MEM_reg_N62) );
  AOI22X1 U4558 ( .A(reg_read_data_1_EX[25]), .B(n3947), .C(alu_result_MEM[25]), .D(n2814), .Y(n3706) );
  OAI21X1 U4559 ( .A(n5189), .B(n3733), .C(n3706), .Y(n4149) );
  OAI21X1 U4560 ( .A(n3720), .B(n3776), .C(n3943), .Y(n3707) );
  AOI21X1 U4561 ( .A(n3941), .B(reg_read_data_2_EX[25]), .C(n3707), .Y(n3708)
         );
  OAI21X1 U4562 ( .A(n5189), .B(n3736), .C(n3708), .Y(n4196) );
  XOR2X1 U4563 ( .A(n4259), .B(n4196), .Y(n3738) );
  AOI22X1 U4564 ( .A(reg_read_data_1_EX[24]), .B(n3947), .C(alu_result_MEM[24]), .D(n2814), .Y(n3709) );
  OAI21X1 U4565 ( .A(n5186), .B(n3733), .C(n3709), .Y(n3993) );
  AOI22X1 U4566 ( .A(alu_result_MEM[24]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[24]), .Y(n3710) );
  AND2X2 U4567 ( .A(n3943), .B(n3710), .Y(n3711) );
  OAI21X1 U4568 ( .A(n5186), .B(n3736), .C(n3711), .Y(n4165) );
  XOR2X1 U4569 ( .A(n4259), .B(n4165), .Y(n3989) );
  FAX1 U4570 ( .A(n4160), .B(n3713), .C(n3712), .YC(n3988), .YS(n3704) );
  NAND2X1 U4571 ( .A(n4149), .B(n4196), .Y(n3715) );
  OAI21X1 U4572 ( .A(n4149), .B(n4196), .C(n3739), .Y(n3714) );
  OAI21X1 U4573 ( .A(n3715), .B(n3953), .C(n3714), .Y(n3716) );
  AOI21X1 U4574 ( .A(n4263), .B(n3717), .C(n3716), .Y(n3718) );
  INVX1 U4575 ( .A(n3718), .Y(inst_EX2MEM_reg_N64) );
  AOI22X1 U4576 ( .A(reg_read_data_1_EX[30]), .B(n3947), .C(alu_result_MEM[30]), .D(n2814), .Y(n3719) );
  OAI21X1 U4577 ( .A(n5231), .B(n2901), .C(n3719), .Y(n4167) );
  OAI21X1 U4578 ( .A(n3720), .B(n3770), .C(n3943), .Y(n3721) );
  AOI21X1 U4579 ( .A(n3941), .B(reg_read_data_2_EX[30]), .C(n3721), .Y(n3722)
         );
  OAI21X1 U4580 ( .A(n5231), .B(n3736), .C(n3722), .Y(n4168) );
  XOR2X1 U4581 ( .A(n4259), .B(n4168), .Y(n3940) );
  AOI22X1 U4582 ( .A(reg_read_data_1_EX[29]), .B(n3947), .C(alu_result_MEM[29]), .D(n2814), .Y(n3723) );
  OAI21X1 U4583 ( .A(n5121), .B(n2901), .C(n3723), .Y(n3963) );
  AOI22X1 U4584 ( .A(alu_result_MEM[29]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[29]), .Y(n3724) );
  OAI21X1 U4585 ( .A(n5121), .B(n3736), .C(n3725), .Y(n4176) );
  XOR2X1 U4586 ( .A(n4259), .B(n4176), .Y(n3959) );
  AOI22X1 U4587 ( .A(reg_read_data_1_EX[28]), .B(n3947), .C(alu_result_MEM[28]), .D(n2814), .Y(n3726) );
  OAI21X1 U4588 ( .A(n5198), .B(n3733), .C(n3726), .Y(n4207) );
  AOI22X1 U4589 ( .A(alu_result_MEM[28]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[28]), .Y(n3727) );
  OAI21X1 U4590 ( .A(n5198), .B(n3736), .C(n3728), .Y(n4150) );
  XOR2X1 U4591 ( .A(n4259), .B(n4150), .Y(n3967) );
  AOI22X1 U4592 ( .A(reg_read_data_1_EX[27]), .B(n3947), .C(alu_result_MEM[27]), .D(n2814), .Y(n3729) );
  OAI21X1 U4593 ( .A(n5195), .B(n2901), .C(n3729), .Y(n4151) );
  AOI22X1 U4594 ( .A(alu_result_MEM[27]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[27]), .Y(n3730) );
  OAI21X1 U4595 ( .A(n5195), .B(n3736), .C(n3731), .Y(n4171) );
  XOR2X1 U4596 ( .A(n4259), .B(n4171), .Y(n3974) );
  AOI22X1 U4597 ( .A(reg_read_data_1_EX[26]), .B(n3947), .C(alu_result_MEM[26]), .D(n2814), .Y(n3732) );
  OAI21X1 U4598 ( .A(n5192), .B(n3733), .C(n3732), .Y(n3985) );
  AOI22X1 U4599 ( .A(n3941), .B(reg_read_data_2_EX[26]), .C(alu_result_MEM[26]), .D(n3942), .Y(n3734) );
  AND2X2 U4600 ( .A(n3943), .B(n3734), .Y(n3735) );
  OAI21X1 U4601 ( .A(n5192), .B(n3736), .C(n3735), .Y(n4173) );
  XOR2X1 U4602 ( .A(n4259), .B(n4173), .Y(n3981) );
  FAX1 U4603 ( .A(n4149), .B(n3738), .C(n3737), .YC(n3980), .YS(n3717) );
  NAND2X1 U4604 ( .A(n4167), .B(n4168), .Y(n3741) );
  OAI21X1 U4605 ( .A(n4167), .B(n4168), .C(n3739), .Y(n3740) );
  OAI21X1 U4606 ( .A(n3741), .B(n4047), .C(n3740), .Y(n3742) );
  AOI21X1 U4607 ( .A(n4263), .B(n3743), .C(n3742), .Y(n3744) );
  INVX1 U4608 ( .A(n3744), .Y(inst_EX2MEM_reg_N69) );
  INVX2 U4609 ( .A(n4426), .Y(n3774) );
  NOR2X1 U4610 ( .A(n3745), .B(n3774), .Y(inst_EX2MEM_reg_N133) );
  NOR2X1 U4611 ( .A(n3746), .B(n2809), .Y(inst_EX2MEM_reg_N132) );
  NOR2X1 U4612 ( .A(n3747), .B(n3774), .Y(inst_EX2MEM_reg_N131) );
  NOR2X1 U4613 ( .A(n3748), .B(n2809), .Y(inst_EX2MEM_reg_N130) );
  NOR2X1 U4614 ( .A(n3749), .B(n3774), .Y(inst_EX2MEM_reg_N129) );
  NOR2X1 U4615 ( .A(n3750), .B(n2809), .Y(inst_EX2MEM_reg_N128) );
  NOR2X1 U4616 ( .A(n3751), .B(n3774), .Y(inst_EX2MEM_reg_N127) );
  NOR2X1 U4617 ( .A(n3752), .B(n2809), .Y(inst_EX2MEM_reg_N126) );
  NOR2X1 U4618 ( .A(n3753), .B(n3774), .Y(inst_EX2MEM_reg_N125) );
  NOR2X1 U4619 ( .A(n3754), .B(n2809), .Y(inst_EX2MEM_reg_N124) );
  NOR2X1 U4620 ( .A(n4419), .B(n3774), .Y(inst_EX2MEM_reg_N123) );
  NOR2X1 U4621 ( .A(n3755), .B(n2809), .Y(inst_EX2MEM_reg_N122) );
  NOR2X1 U4622 ( .A(n3756), .B(n3774), .Y(inst_EX2MEM_reg_N121) );
  NOR2X1 U4623 ( .A(n4375), .B(n2809), .Y(inst_EX2MEM_reg_N120) );
  NOR2X1 U4624 ( .A(n3757), .B(n3774), .Y(inst_EX2MEM_reg_N119) );
  NOR2X1 U4625 ( .A(n3758), .B(n3774), .Y(inst_EX2MEM_reg_N118) );
  NOR2X1 U4626 ( .A(n4367), .B(n2809), .Y(inst_EX2MEM_reg_N117) );
  NOR2X1 U4627 ( .A(n3759), .B(n3774), .Y(inst_EX2MEM_reg_N116) );
  NOR2X1 U4628 ( .A(n3760), .B(n2809), .Y(inst_EX2MEM_reg_N115) );
  NOR2X1 U4629 ( .A(n3761), .B(n3774), .Y(inst_EX2MEM_reg_N114) );
  NOR2X1 U4630 ( .A(n3762), .B(n2809), .Y(inst_EX2MEM_reg_N113) );
  NOR2X1 U4631 ( .A(n3763), .B(n3774), .Y(inst_EX2MEM_reg_N112) );
  NOR2X1 U4632 ( .A(n3764), .B(n2809), .Y(inst_EX2MEM_reg_N111) );
  NOR2X1 U4633 ( .A(n3765), .B(n3774), .Y(inst_EX2MEM_reg_N110) );
  NOR2X1 U4634 ( .A(n3766), .B(n2809), .Y(inst_EX2MEM_reg_N109) );
  NOR2X1 U4635 ( .A(n4332), .B(n3774), .Y(inst_EX2MEM_reg_N108) );
  NOR2X1 U4636 ( .A(n3767), .B(n3774), .Y(u_MEM2WB_reg_N6) );
  NOR2X1 U4637 ( .A(n4429), .B(n2809), .Y(u_MEM2WB_reg_N5) );
  NOR2X1 U4638 ( .A(n3768), .B(n3805), .Y(u_MEM2WB_reg_N4) );
  NOR2X1 U4639 ( .A(n4430), .B(n3774), .Y(u_MEM2WB_reg_N3) );
  NOR2X1 U4640 ( .A(n3769), .B(n2809), .Y(u_MEM2WB_reg_N70) );
  NOR2X1 U4641 ( .A(n3770), .B(n3774), .Y(u_MEM2WB_reg_N69) );
  NOR2X1 U4642 ( .A(n3771), .B(n3805), .Y(u_MEM2WB_reg_N68) );
  NOR2X1 U4643 ( .A(n3772), .B(n2809), .Y(u_MEM2WB_reg_N67) );
  NOR2X1 U4644 ( .A(n3773), .B(n3774), .Y(u_MEM2WB_reg_N66) );
  INVX1 U4645 ( .A(alu_result_MEM[26]), .Y(n3775) );
  NOR2X1 U4646 ( .A(n3775), .B(n2809), .Y(u_MEM2WB_reg_N65) );
  NOR2X1 U4647 ( .A(n3776), .B(n2809), .Y(u_MEM2WB_reg_N64) );
  NOR2X1 U4648 ( .A(n3777), .B(n2809), .Y(u_MEM2WB_reg_N63) );
  NOR2X1 U4649 ( .A(n3778), .B(n2809), .Y(u_MEM2WB_reg_N62) );
  NOR2X1 U4650 ( .A(n3779), .B(n2809), .Y(u_MEM2WB_reg_N61) );
  NOR2X1 U4651 ( .A(n3780), .B(n2809), .Y(u_MEM2WB_reg_N60) );
  NOR2X1 U4652 ( .A(n3781), .B(n2809), .Y(u_MEM2WB_reg_N59) );
  INVX1 U4653 ( .A(alu_result_MEM[19]), .Y(n3782) );
  NOR2X1 U4654 ( .A(n3782), .B(n2809), .Y(u_MEM2WB_reg_N58) );
  NOR2X1 U4655 ( .A(n3783), .B(n2809), .Y(u_MEM2WB_reg_N57) );
  NOR2X1 U4656 ( .A(n3784), .B(n3774), .Y(u_MEM2WB_reg_N56) );
  NOR2X1 U4657 ( .A(n3785), .B(n2809), .Y(u_MEM2WB_reg_N55) );
  NOR2X1 U4658 ( .A(n3786), .B(n3774), .Y(u_MEM2WB_reg_N54) );
  NOR2X1 U4659 ( .A(n3787), .B(n2809), .Y(u_MEM2WB_reg_N53) );
  NOR2X1 U4660 ( .A(n3788), .B(n3774), .Y(u_MEM2WB_reg_N52) );
  NOR2X1 U4661 ( .A(n3789), .B(n2809), .Y(u_MEM2WB_reg_N51) );
  NOR2X1 U4662 ( .A(n3790), .B(n3774), .Y(u_MEM2WB_reg_N50) );
  NOR2X1 U4663 ( .A(n3791), .B(n3774), .Y(u_MEM2WB_reg_N49) );
  NOR2X1 U4664 ( .A(n3792), .B(n2809), .Y(u_MEM2WB_reg_N48) );
  NOR2X1 U4665 ( .A(n3793), .B(n3774), .Y(u_MEM2WB_reg_N47) );
  NOR2X1 U4666 ( .A(n3794), .B(n2809), .Y(u_MEM2WB_reg_N46) );
  NOR2X1 U4667 ( .A(n3795), .B(n3774), .Y(u_MEM2WB_reg_N45) );
  INVX1 U4668 ( .A(alu_result_MEM[5]), .Y(n3796) );
  NOR2X1 U4669 ( .A(n3796), .B(n3774), .Y(u_MEM2WB_reg_N44) );
  NOR2X1 U4670 ( .A(n3797), .B(n2809), .Y(u_MEM2WB_reg_N43) );
  NOR2X1 U4671 ( .A(n3798), .B(n3774), .Y(u_MEM2WB_reg_N42) );
  NOR2X1 U4672 ( .A(n4432), .B(n3774), .Y(u_MEM2WB_reg_N41) );
  NOR2X1 U4673 ( .A(n4434), .B(n2809), .Y(u_MEM2WB_reg_N40) );
  NOR2X1 U4674 ( .A(n4443), .B(n3774), .Y(u_MEM2WB_reg_N39) );
  INVX1 U4675 ( .A(reg_write_address_MEM[4]), .Y(n3799) );
  NOR2X1 U4676 ( .A(n3799), .B(n2809), .Y(u_MEM2WB_reg_N75) );
  NOR2X1 U4677 ( .A(n3800), .B(n3774), .Y(u_MEM2WB_reg_N74) );
  NOR2X1 U4678 ( .A(n3801), .B(n3774), .Y(u_MEM2WB_reg_N73) );
  NOR2X1 U4679 ( .A(n3802), .B(n2809), .Y(u_MEM2WB_reg_N72) );
  NOR2X1 U4680 ( .A(n3803), .B(n3774), .Y(u_MEM2WB_reg_N71) );
  NOR2X1 U4681 ( .A(n3804), .B(n2809), .Y(inst_EX2MEM_reg_N6) );
  INVX1 U4682 ( .A(op_type_EX[0]), .Y(n4192) );
  NOR2X1 U4683 ( .A(n4192), .B(n2809), .Y(inst_EX2MEM_reg_N3) );
  INVX1 U4684 ( .A(reg_read_data_2_EX[31]), .Y(n3806) );
  NOR2X1 U4685 ( .A(n3806), .B(n2809), .Y(inst_EX2MEM_reg_N102) );
  INVX1 U4686 ( .A(reg_read_data_2_EX[30]), .Y(n3807) );
  NOR2X1 U4687 ( .A(n3807), .B(n3805), .Y(inst_EX2MEM_reg_N101) );
  INVX1 U4688 ( .A(reg_read_data_2_EX[29]), .Y(n3808) );
  NOR2X1 U4689 ( .A(n3808), .B(n2809), .Y(inst_EX2MEM_reg_N100) );
  INVX1 U4690 ( .A(reg_read_data_2_EX[28]), .Y(n3809) );
  NOR2X1 U4691 ( .A(n3809), .B(n3805), .Y(inst_EX2MEM_reg_N99) );
  INVX1 U4692 ( .A(reg_read_data_2_EX[27]), .Y(n3810) );
  NOR2X1 U4693 ( .A(n3810), .B(n3805), .Y(inst_EX2MEM_reg_N98) );
  INVX1 U4694 ( .A(reg_read_data_2_EX[26]), .Y(n3811) );
  NOR2X1 U4695 ( .A(n3811), .B(n2809), .Y(inst_EX2MEM_reg_N97) );
  INVX1 U4696 ( .A(reg_read_data_2_EX[25]), .Y(n3812) );
  NOR2X1 U4697 ( .A(n3812), .B(n2809), .Y(inst_EX2MEM_reg_N96) );
  INVX1 U4698 ( .A(reg_read_data_2_EX[24]), .Y(n3813) );
  NOR2X1 U4699 ( .A(n3813), .B(n3805), .Y(inst_EX2MEM_reg_N95) );
  INVX1 U4700 ( .A(reg_read_data_2_EX[23]), .Y(n3814) );
  NOR2X1 U4701 ( .A(n3814), .B(n2809), .Y(inst_EX2MEM_reg_N94) );
  INVX1 U4702 ( .A(reg_read_data_2_EX[22]), .Y(n3815) );
  NOR2X1 U4703 ( .A(n3815), .B(n3805), .Y(inst_EX2MEM_reg_N93) );
  INVX1 U4704 ( .A(reg_read_data_2_EX[21]), .Y(n3816) );
  NOR2X1 U4705 ( .A(n3816), .B(n3805), .Y(inst_EX2MEM_reg_N92) );
  INVX1 U4706 ( .A(reg_read_data_2_EX[20]), .Y(n3817) );
  NOR2X1 U4707 ( .A(n3817), .B(n3805), .Y(inst_EX2MEM_reg_N91) );
  INVX1 U4708 ( .A(reg_read_data_2_EX[19]), .Y(n3818) );
  NOR2X1 U4709 ( .A(n3818), .B(n3805), .Y(inst_EX2MEM_reg_N90) );
  INVX1 U4710 ( .A(reg_read_data_2_EX[18]), .Y(n3819) );
  NOR2X1 U4711 ( .A(n3819), .B(n3805), .Y(inst_EX2MEM_reg_N89) );
  INVX1 U4712 ( .A(reg_read_data_2_EX[17]), .Y(n3820) );
  NOR2X1 U4713 ( .A(n3820), .B(n3805), .Y(inst_EX2MEM_reg_N88) );
  INVX1 U4714 ( .A(reg_read_data_2_EX[16]), .Y(n3821) );
  NOR2X1 U4715 ( .A(n3821), .B(n3805), .Y(inst_EX2MEM_reg_N87) );
  INVX1 U4716 ( .A(reg_read_data_2_EX[15]), .Y(n3822) );
  NOR2X1 U4717 ( .A(n3822), .B(n3805), .Y(inst_EX2MEM_reg_N86) );
  INVX1 U4718 ( .A(reg_read_data_2_EX[14]), .Y(n3823) );
  NOR2X1 U4719 ( .A(n3823), .B(n3805), .Y(inst_EX2MEM_reg_N85) );
  INVX1 U4720 ( .A(reg_read_data_2_EX[13]), .Y(n3824) );
  NOR2X1 U4721 ( .A(n3824), .B(n3805), .Y(inst_EX2MEM_reg_N84) );
  INVX1 U4722 ( .A(reg_read_data_2_EX[12]), .Y(n3825) );
  NOR2X1 U4723 ( .A(n3825), .B(n3805), .Y(inst_EX2MEM_reg_N83) );
  INVX1 U4724 ( .A(reg_read_data_2_EX[11]), .Y(n3826) );
  NOR2X1 U4725 ( .A(n3826), .B(n3805), .Y(inst_EX2MEM_reg_N82) );
  INVX1 U4726 ( .A(reg_read_data_2_EX[10]), .Y(n3827) );
  NOR2X1 U4727 ( .A(n3827), .B(n3805), .Y(inst_EX2MEM_reg_N81) );
  INVX1 U4728 ( .A(reg_read_data_2_EX[9]), .Y(n3828) );
  NOR2X1 U4729 ( .A(n3828), .B(n3805), .Y(inst_EX2MEM_reg_N80) );
  INVX1 U4730 ( .A(reg_read_data_2_EX[8]), .Y(n3829) );
  NOR2X1 U4731 ( .A(n3829), .B(n3805), .Y(inst_EX2MEM_reg_N79) );
  INVX1 U4732 ( .A(reg_read_data_2_EX[7]), .Y(n3830) );
  NOR2X1 U4733 ( .A(n3830), .B(n3805), .Y(inst_EX2MEM_reg_N78) );
  INVX1 U4734 ( .A(reg_read_data_2_EX[6]), .Y(n3831) );
  NOR2X1 U4735 ( .A(n3831), .B(n2809), .Y(inst_EX2MEM_reg_N77) );
  INVX1 U4736 ( .A(reg_read_data_2_EX[5]), .Y(n3832) );
  NOR2X1 U4737 ( .A(n3832), .B(n3805), .Y(inst_EX2MEM_reg_N76) );
  INVX1 U4738 ( .A(reg_read_data_2_EX[4]), .Y(n3833) );
  NOR2X1 U4739 ( .A(n3833), .B(n2809), .Y(inst_EX2MEM_reg_N75) );
  INVX1 U4740 ( .A(reg_read_data_2_EX[3]), .Y(n3834) );
  NOR2X1 U4741 ( .A(n3834), .B(n3805), .Y(inst_EX2MEM_reg_N74) );
  INVX1 U4742 ( .A(reg_read_data_2_EX[2]), .Y(n3835) );
  NOR2X1 U4743 ( .A(n3835), .B(n2809), .Y(inst_EX2MEM_reg_N73) );
  INVX1 U4744 ( .A(reg_read_data_2_EX[1]), .Y(n3836) );
  NOR2X1 U4745 ( .A(n3836), .B(n3805), .Y(inst_EX2MEM_reg_N72) );
  INVX1 U4746 ( .A(reg_read_data_2_EX[0]), .Y(n3837) );
  NOR2X1 U4747 ( .A(n3837), .B(n2809), .Y(inst_EX2MEM_reg_N71) );
  NOR2X1 U4748 ( .A(n3838), .B(n3805), .Y(inst_EX2MEM_reg_N107) );
  NOR2X1 U4749 ( .A(n3839), .B(n2809), .Y(inst_EX2MEM_reg_N106) );
  NOR2X1 U4750 ( .A(n3840), .B(n3805), .Y(inst_EX2MEM_reg_N105) );
  NOR2X1 U4751 ( .A(n3841), .B(n2809), .Y(inst_EX2MEM_reg_N104) );
  NOR2X1 U4752 ( .A(n3842), .B(n3805), .Y(inst_EX2MEM_reg_N103) );
  INVX1 U4753 ( .A(instruction_ID[5]), .Y(n4672) );
  NOR2X1 U4754 ( .A(n4312), .B(n4672), .Y(inst_ID2EX_reg_N108) );
  INVX1 U4755 ( .A(inst_addr_ID[31]), .Y(n4683) );
  NOR2X1 U4756 ( .A(n4312), .B(n4683), .Y(inst_ID2EX_reg_N38) );
  INVX1 U4757 ( .A(inst_addr_ID[30]), .Y(n4685) );
  NOR2X1 U4758 ( .A(n4312), .B(n4685), .Y(inst_ID2EX_reg_N37) );
  INVX1 U4759 ( .A(inst_addr_ID[29]), .Y(n4689) );
  NOR2X1 U4760 ( .A(n4312), .B(n4689), .Y(inst_ID2EX_reg_N36) );
  INVX1 U4761 ( .A(inst_addr_ID[28]), .Y(n4690) );
  NOR2X1 U4762 ( .A(n4312), .B(n4690), .Y(inst_ID2EX_reg_N35) );
  INVX1 U4763 ( .A(inst_addr_ID[27]), .Y(n4692) );
  NOR2X1 U4764 ( .A(n3844), .B(n4692), .Y(inst_ID2EX_reg_N34) );
  INVX1 U4765 ( .A(inst_addr_ID[26]), .Y(n4693) );
  NOR2X1 U4766 ( .A(n3844), .B(n4693), .Y(inst_ID2EX_reg_N33) );
  INVX1 U4767 ( .A(inst_addr_ID[25]), .Y(n4695) );
  NOR2X1 U4768 ( .A(n3844), .B(n4695), .Y(inst_ID2EX_reg_N32) );
  INVX1 U4769 ( .A(inst_addr_ID[24]), .Y(n4697) );
  NOR2X1 U4770 ( .A(n3844), .B(n4697), .Y(inst_ID2EX_reg_N31) );
  INVX1 U4771 ( .A(inst_addr_ID[23]), .Y(n4699) );
  NOR2X1 U4772 ( .A(n3844), .B(n4699), .Y(inst_ID2EX_reg_N30) );
  INVX1 U4773 ( .A(inst_addr_ID[22]), .Y(n4701) );
  NOR2X1 U4774 ( .A(n3844), .B(n4701), .Y(inst_ID2EX_reg_N29) );
  INVX1 U4775 ( .A(inst_addr_ID[21]), .Y(n4703) );
  NOR2X1 U4776 ( .A(n3844), .B(n4703), .Y(inst_ID2EX_reg_N28) );
  INVX1 U4777 ( .A(inst_addr_ID[20]), .Y(n4706) );
  NOR2X1 U4778 ( .A(n3844), .B(n4706), .Y(inst_ID2EX_reg_N27) );
  INVX1 U4779 ( .A(inst_addr_ID[19]), .Y(n4708) );
  NOR2X1 U4780 ( .A(n3844), .B(n4708), .Y(inst_ID2EX_reg_N26) );
  INVX1 U4781 ( .A(inst_addr_ID[18]), .Y(n4710) );
  NOR2X1 U4782 ( .A(n3844), .B(n4710), .Y(inst_ID2EX_reg_N25) );
  INVX1 U4783 ( .A(inst_addr_ID[17]), .Y(n4712) );
  NOR2X1 U4784 ( .A(n3844), .B(n4712), .Y(inst_ID2EX_reg_N24) );
  INVX1 U4785 ( .A(inst_addr_ID[16]), .Y(n4714) );
  NOR2X1 U4786 ( .A(n3844), .B(n4714), .Y(inst_ID2EX_reg_N23) );
  INVX1 U4787 ( .A(inst_addr_ID[15]), .Y(n4716) );
  NOR2X1 U4788 ( .A(n3843), .B(n4716), .Y(inst_ID2EX_reg_N22) );
  INVX1 U4789 ( .A(inst_addr_ID[14]), .Y(n4718) );
  NOR2X1 U4790 ( .A(n3843), .B(n4718), .Y(inst_ID2EX_reg_N21) );
  INVX1 U4791 ( .A(inst_addr_ID[13]), .Y(n4720) );
  NOR2X1 U4792 ( .A(n3843), .B(n4720), .Y(inst_ID2EX_reg_N20) );
  INVX1 U4793 ( .A(inst_addr_ID[12]), .Y(n4722) );
  NOR2X1 U4794 ( .A(n3843), .B(n4722), .Y(inst_ID2EX_reg_N19) );
  INVX1 U4795 ( .A(inst_addr_ID[11]), .Y(n4724) );
  NOR2X1 U4796 ( .A(n3843), .B(n4724), .Y(inst_ID2EX_reg_N18) );
  INVX1 U4797 ( .A(inst_addr_ID[10]), .Y(n4726) );
  NOR2X1 U4798 ( .A(n3843), .B(n4726), .Y(inst_ID2EX_reg_N17) );
  INVX1 U4799 ( .A(inst_addr_ID[9]), .Y(n4729) );
  NOR2X1 U4800 ( .A(n3843), .B(n4729), .Y(inst_ID2EX_reg_N16) );
  INVX1 U4801 ( .A(inst_addr_ID[8]), .Y(n4731) );
  NOR2X1 U4802 ( .A(n3843), .B(n4731), .Y(inst_ID2EX_reg_N15) );
  INVX1 U4803 ( .A(inst_addr_ID[7]), .Y(n4733) );
  NOR2X1 U4804 ( .A(n3843), .B(n4733), .Y(inst_ID2EX_reg_N14) );
  INVX1 U4805 ( .A(inst_addr_ID[6]), .Y(n4735) );
  NOR2X1 U4806 ( .A(n3843), .B(n4735), .Y(inst_ID2EX_reg_N13) );
  INVX1 U4807 ( .A(inst_addr_ID[5]), .Y(n4737) );
  NOR2X1 U4808 ( .A(n3843), .B(n4737), .Y(inst_ID2EX_reg_N12) );
  INVX1 U4809 ( .A(inst_addr_ID[4]), .Y(n4739) );
  NOR2X1 U4810 ( .A(n3843), .B(n4739), .Y(inst_ID2EX_reg_N11) );
  INVX1 U4811 ( .A(inst_addr_ID[3]), .Y(n4741) );
  NOR2X1 U4812 ( .A(n3843), .B(n4741), .Y(inst_ID2EX_reg_N10) );
  INVX1 U4813 ( .A(inst_addr_ID[2]), .Y(n4743) );
  NOR2X1 U4814 ( .A(n3845), .B(n4743), .Y(inst_ID2EX_reg_N9) );
  INVX1 U4815 ( .A(inst_addr_ID[1]), .Y(n4744) );
  NOR2X1 U4816 ( .A(n3845), .B(n4744), .Y(inst_ID2EX_reg_N8) );
  INVX1 U4817 ( .A(inst_addr_ID[0]), .Y(n4746) );
  NOR2X1 U4818 ( .A(n3845), .B(n4746), .Y(inst_ID2EX_reg_N7) );
  INVX1 U4819 ( .A(instruction_ID[15]), .Y(n4652) );
  NOR2X1 U4820 ( .A(n3845), .B(n4652), .Y(inst_ID2EX_reg_N134) );
  INVX1 U4821 ( .A(instruction_ID[14]), .Y(n4654) );
  NOR2X1 U4822 ( .A(n3845), .B(n4654), .Y(inst_ID2EX_reg_N117) );
  INVX1 U4823 ( .A(instruction_ID[13]), .Y(n4656) );
  NOR2X1 U4824 ( .A(n3844), .B(n4656), .Y(inst_ID2EX_reg_N116) );
  INVX1 U4825 ( .A(instruction_ID[12]), .Y(n4658) );
  NOR2X1 U4826 ( .A(n3845), .B(n4658), .Y(inst_ID2EX_reg_N115) );
  INVX1 U4827 ( .A(instruction_ID[11]), .Y(n4660) );
  NOR2X1 U4828 ( .A(n3843), .B(n4660), .Y(inst_ID2EX_reg_N114) );
  INVX1 U4829 ( .A(instruction_ID[10]), .Y(n4662) );
  NOR2X1 U4830 ( .A(n3844), .B(n4662), .Y(inst_ID2EX_reg_N113) );
  INVX1 U4831 ( .A(instruction_ID[9]), .Y(n4664) );
  NOR2X1 U4832 ( .A(n3845), .B(n4664), .Y(inst_ID2EX_reg_N112) );
  INVX1 U4833 ( .A(instruction_ID[8]), .Y(n4666) );
  NOR2X1 U4834 ( .A(n3843), .B(n4666), .Y(inst_ID2EX_reg_N111) );
  INVX1 U4835 ( .A(instruction_ID[7]), .Y(n4668) );
  NOR2X1 U4836 ( .A(n3844), .B(n4668), .Y(inst_ID2EX_reg_N110) );
  INVX1 U4837 ( .A(instruction_ID[6]), .Y(n4670) );
  NOR2X1 U4838 ( .A(n3845), .B(n4670), .Y(inst_ID2EX_reg_N109) );
  INVX1 U4839 ( .A(instruction_ID[4]), .Y(n4674) );
  NOR2X1 U4840 ( .A(n3845), .B(n4674), .Y(inst_ID2EX_reg_N107) );
  INVX1 U4841 ( .A(n2795), .Y(n3845) );
  INVX1 U4842 ( .A(instruction_ID[3]), .Y(n4676) );
  NOR2X1 U4843 ( .A(n3845), .B(n4676), .Y(inst_ID2EX_reg_N106) );
  INVX1 U4844 ( .A(instruction_ID[2]), .Y(n4678) );
  NOR2X1 U4845 ( .A(n3845), .B(n4678), .Y(inst_ID2EX_reg_N105) );
  INVX1 U4846 ( .A(instruction_ID[1]), .Y(n4680) );
  NOR2X1 U4847 ( .A(n3845), .B(n4680), .Y(inst_ID2EX_reg_N104) );
  INVX1 U4848 ( .A(instruction_ID[0]), .Y(n4682) );
  NOR2X1 U4849 ( .A(n4312), .B(n4682), .Y(inst_ID2EX_reg_N103) );
  NOR2X1 U4850 ( .A(n4642), .B(n5524), .Y(inst_ID2EX_reg_N139) );
  NOR2X1 U4851 ( .A(n4644), .B(n5524), .Y(inst_ID2EX_reg_N138) );
  NOR2X1 U4852 ( .A(n4646), .B(n5524), .Y(inst_ID2EX_reg_N137) );
  NOR2X1 U4853 ( .A(n4648), .B(n5524), .Y(inst_ID2EX_reg_N136) );
  NOR2X1 U4854 ( .A(n4650), .B(n5524), .Y(inst_ID2EX_reg_N135) );
  NOR2X1 U4855 ( .A(n4632), .B(n5524), .Y(inst_ID2EX_reg_N170) );
  NOR2X1 U4856 ( .A(n4634), .B(n5524), .Y(inst_ID2EX_reg_N169) );
  NOR2X1 U4857 ( .A(n4636), .B(n5524), .Y(inst_ID2EX_reg_N168) );
  NOR2X1 U4858 ( .A(n4638), .B(n5524), .Y(inst_ID2EX_reg_N167) );
  NOR2X1 U4859 ( .A(n4640), .B(n5524), .Y(inst_ID2EX_reg_N166) );
  NOR2X1 U4860 ( .A(inst_address[24]), .B(n5524), .Y(n3858) );
  NOR2X1 U4861 ( .A(inst_address[22]), .B(n5524), .Y(n3857) );
  NOR2X1 U4862 ( .A(inst_address[20]), .B(n5524), .Y(n3856) );
  NOR2X1 U4863 ( .A(inst_address[18]), .B(n5524), .Y(n3855) );
  NOR2X1 U4864 ( .A(n3846), .B(n4719), .Y(n3852) );
  NOR2X1 U4865 ( .A(n3847), .B(n4286), .Y(n3849) );
  NAND2X1 U4866 ( .A(inst_address[15]), .B(n3849), .Y(n3848) );
  NOR2X1 U4867 ( .A(inst_address[16]), .B(n3848), .Y(n3904) );
  NOR2X1 U4868 ( .A(n3851), .B(n3850), .Y(n4296) );
  OAI21X1 U4869 ( .A(inst_address[15]), .B(n4299), .C(n4296), .Y(n3903) );
  NOR2X1 U4870 ( .A(n3904), .B(n3903), .Y(n4301) );
  NAND3X1 U4871 ( .A(n3852), .B(inst_address[16]), .C(inst_address[15]), .Y(
        n3853) );
  NOR2X1 U4872 ( .A(n3854), .B(n3853), .Y(n3859) );
  INVX1 U4873 ( .A(inst_address[17]), .Y(n4713) );
  NAND3X1 U4874 ( .A(n3859), .B(n2795), .C(n4713), .Y(n4300) );
  NAND2X1 U4875 ( .A(n4301), .B(n4300), .Y(n3899) );
  NOR2X1 U4876 ( .A(n3855), .B(n3899), .Y(n3891) );
  OAI21X1 U4877 ( .A(inst_address[19]), .B(n5524), .C(n3891), .Y(n3888) );
  NOR2X1 U4878 ( .A(n3856), .B(n3888), .Y(n3880) );
  OAI21X1 U4879 ( .A(inst_address[21]), .B(n3933), .C(n3880), .Y(n3877) );
  NOR2X1 U4880 ( .A(n3857), .B(n3877), .Y(n3869) );
  OAI21X1 U4881 ( .A(inst_address[23]), .B(n5524), .C(n3869), .Y(n3866) );
  NOR2X1 U4882 ( .A(n3858), .B(n3866), .Y(n5503) );
  INVX1 U4883 ( .A(n5503), .Y(n3861) );
  NOR2X1 U4884 ( .A(inst_address[25]), .B(n5524), .Y(n3860) );
  INVX1 U4885 ( .A(inst_address[24]), .Y(n4698) );
  INVX1 U4886 ( .A(inst_address[22]), .Y(n4702) );
  INVX1 U4887 ( .A(inst_address[20]), .Y(n4707) );
  INVX1 U4888 ( .A(inst_address[18]), .Y(n4711) );
  NAND2X1 U4889 ( .A(n3859), .B(inst_address[17]), .Y(n3897) );
  NOR2X1 U4890 ( .A(n4711), .B(n3897), .Y(n3892) );
  NAND2X1 U4891 ( .A(inst_address[19]), .B(n3892), .Y(n3886) );
  NOR2X1 U4892 ( .A(n4707), .B(n3886), .Y(n3881) );
  NAND2X1 U4893 ( .A(inst_address[21]), .B(n3881), .Y(n3875) );
  NOR2X1 U4894 ( .A(n4702), .B(n3875), .Y(n3870) );
  NAND2X1 U4895 ( .A(inst_address[23]), .B(n3870), .Y(n3864) );
  NOR2X1 U4896 ( .A(n4698), .B(n3864), .Y(n4615) );
  AOI22X1 U4897 ( .A(inst_address[25]), .B(n3861), .C(n3860), .D(n4615), .Y(
        n3863) );
  AOI22X1 U4898 ( .A(n4294), .B(shifted_address_MEM[25]), .C(n3902), .D(
        jump_inst_addr_MEM[25]), .Y(n3862) );
  NAND2X1 U4899 ( .A(n3863), .B(n3862), .Y(n2189) );
  OAI21X1 U4900 ( .A(n3933), .B(n3864), .C(n4698), .Y(n3865) );
  OAI21X1 U4901 ( .A(n4698), .B(n3866), .C(n3865), .Y(n3868) );
  AOI22X1 U4902 ( .A(n4294), .B(shifted_address_MEM[24]), .C(n3902), .D(
        jump_inst_addr_MEM[24]), .Y(n3867) );
  NAND2X1 U4903 ( .A(n3868), .B(n3867), .Y(n2190) );
  INVX1 U4904 ( .A(n3869), .Y(n3872) );
  NOR2X1 U4905 ( .A(inst_address[23]), .B(n3933), .Y(n3871) );
  AOI22X1 U4906 ( .A(inst_address[23]), .B(n3872), .C(n3871), .D(n3870), .Y(
        n3874) );
  AOI22X1 U4907 ( .A(n4294), .B(shifted_address_MEM[23]), .C(n3902), .D(
        jump_inst_addr_MEM[23]), .Y(n3873) );
  NAND2X1 U4908 ( .A(n3874), .B(n3873), .Y(n2191) );
  OAI21X1 U4909 ( .A(n3933), .B(n3875), .C(n4702), .Y(n3876) );
  OAI21X1 U4910 ( .A(n4702), .B(n3877), .C(n3876), .Y(n3879) );
  AOI22X1 U4911 ( .A(n4294), .B(shifted_address_MEM[22]), .C(n3902), .D(
        jump_inst_addr_MEM[22]), .Y(n3878) );
  NAND2X1 U4912 ( .A(n3879), .B(n3878), .Y(n2192) );
  INVX1 U4913 ( .A(n3880), .Y(n3883) );
  NOR2X1 U4914 ( .A(inst_address[21]), .B(n3933), .Y(n3882) );
  AOI22X1 U4915 ( .A(inst_address[21]), .B(n3883), .C(n3882), .D(n3881), .Y(
        n3885) );
  AOI22X1 U4916 ( .A(n4294), .B(shifted_address_MEM[21]), .C(n3902), .D(
        jump_inst_addr_MEM[21]), .Y(n3884) );
  NAND2X1 U4917 ( .A(n3885), .B(n3884), .Y(n2193) );
  OAI21X1 U4918 ( .A(n4312), .B(n3886), .C(n4707), .Y(n3887) );
  OAI21X1 U4919 ( .A(n4707), .B(n3888), .C(n3887), .Y(n3890) );
  AOI22X1 U4920 ( .A(n4294), .B(shifted_address_MEM[20]), .C(n3902), .D(
        jump_inst_addr_MEM[20]), .Y(n3889) );
  NAND2X1 U4921 ( .A(n3890), .B(n3889), .Y(n2194) );
  INVX1 U4922 ( .A(n3891), .Y(n3894) );
  NOR2X1 U4923 ( .A(inst_address[19]), .B(n3933), .Y(n3893) );
  AOI22X1 U4924 ( .A(inst_address[19]), .B(n3894), .C(n3893), .D(n3892), .Y(
        n3896) );
  AOI22X1 U4925 ( .A(n4294), .B(shifted_address_MEM[19]), .C(n3902), .D(
        jump_inst_addr_MEM[19]), .Y(n3895) );
  NAND2X1 U4926 ( .A(n3896), .B(n3895), .Y(n2195) );
  OAI21X1 U4927 ( .A(n4312), .B(n3897), .C(n4711), .Y(n3898) );
  OAI21X1 U4928 ( .A(n4711), .B(n3899), .C(n3898), .Y(n3901) );
  AOI22X1 U4929 ( .A(n4294), .B(shifted_address_MEM[18]), .C(n3902), .D(
        jump_inst_addr_MEM[18]), .Y(n3900) );
  NAND2X1 U4930 ( .A(n3901), .B(n3900), .Y(n2196) );
  AOI22X1 U4931 ( .A(inst_address[16]), .B(n3903), .C(n3902), .D(
        jump_inst_addr_MEM[16]), .Y(n3906) );
  AOI21X1 U4932 ( .A(n5526), .B(shifted_address_MEM[16]), .C(n3904), .Y(n3905)
         );
  NAND2X1 U4933 ( .A(n3906), .B(n3905), .Y(n2198) );
  AOI22X1 U4934 ( .A(n3909), .B(n3908), .C(inst_address[11]), .D(n3907), .Y(
        n3911) );
  AOI22X1 U4935 ( .A(n4294), .B(shifted_address_MEM[11]), .C(n5497), .D(
        jump_inst_addr_MEM[11]), .Y(n3910) );
  NAND2X1 U4936 ( .A(n3911), .B(n3910), .Y(n2203) );
  AOI22X1 U4937 ( .A(n4294), .B(shifted_address_MEM[10]), .C(n5497), .D(
        jump_inst_addr_MEM[10]), .Y(n3916) );
  INVX1 U4938 ( .A(n3913), .Y(n3912) );
  OAI21X1 U4939 ( .A(n3912), .B(n3933), .C(n4727), .Y(n3920) );
  OAI21X1 U4940 ( .A(n4312), .B(n3913), .C(n4728), .Y(n3914) );
  OAI21X1 U4941 ( .A(n4728), .B(n3920), .C(n3914), .Y(n3915) );
  NAND2X1 U4942 ( .A(n3916), .B(n3915), .Y(n2204) );
  AOI22X1 U4943 ( .A(n4294), .B(shifted_address_MEM[9]), .C(n5497), .D(
        jump_inst_addr_MEM[9]), .Y(n3923) );
  INVX1 U4945 ( .A(inst_address[8]), .Y(n4732) );
  NAND2X1 U4946 ( .A(n2795), .B(n3917), .Y(n3928) );
  NOR2X1 U4947 ( .A(n4734), .B(n3928), .Y(n3925) );
  INVX1 U4948 ( .A(inst_address[9]), .Y(n4730) );
  OAI21X1 U4949 ( .A(n4732), .B(n3918), .C(n4730), .Y(n3919) );
  OAI21X1 U4950 ( .A(1'b0), .B(n3920), .C(n3919), .Y(n3922) );
  NAND2X1 U4951 ( .A(n3923), .B(n3922), .Y(n2205) );
  AOI22X1 U4952 ( .A(n4294), .B(shifted_address_MEM[8]), .C(n5497), .D(
        jump_inst_addr_MEM[8]), .Y(n3927) );
  OAI21X1 U4953 ( .A(n3924), .B(n3933), .C(n4727), .Y(n3929) );
  AOI22X1 U4954 ( .A(inst_address[8]), .B(n3929), .C(n3925), .D(n4732), .Y(
        n3926) );
  NAND2X1 U4955 ( .A(n3927), .B(n3926), .Y(n2206) );
  AOI22X1 U4956 ( .A(n4294), .B(shifted_address_MEM[7]), .C(n5497), .D(
        jump_inst_addr_MEM[7]), .Y(n3932) );
  OAI21X1 U4957 ( .A(inst_address[7]), .B(n3930), .C(n3929), .Y(n3931) );
  NAND2X1 U4958 ( .A(n3932), .B(n3931), .Y(n2207) );
  AOI22X1 U4959 ( .A(n4294), .B(shifted_address_MEM[4]), .C(n5497), .D(
        jump_inst_addr_MEM[4]), .Y(n3938) );
  INVX1 U4960 ( .A(inst_address[4]), .Y(n4740) );
  OAI21X1 U4961 ( .A(n3934), .B(n3933), .C(n4727), .Y(n4270) );
  INVX1 U4962 ( .A(n3934), .Y(n3935) );
  OAI21X1 U4963 ( .A(n4312), .B(n3935), .C(n4740), .Y(n3936) );
  OAI21X1 U4964 ( .A(n4740), .B(n4270), .C(n3936), .Y(n3937) );
  NAND2X1 U4965 ( .A(n3938), .B(n3937), .Y(n2210) );
  FAX1 U4966 ( .A(n4167), .B(n3940), .C(n3939), .YC(n3952), .YS(n3743) );
  AOI22X1 U4967 ( .A(alu_result_MEM[31]), .B(n3942), .C(n3941), .D(
        reg_read_data_2_EX[31]), .Y(n3944) );
  NAND2X1 U4968 ( .A(n3944), .B(n3943), .Y(n3945) );
  AOI21X1 U4969 ( .A(n5204), .B(n3946), .C(n3945), .Y(n4190) );
  XOR2X1 U4970 ( .A(n4259), .B(n4162), .Y(n3950) );
  AOI22X1 U4971 ( .A(reg_read_data_1_EX[31]), .B(n3947), .C(alu_result_MEM[31]), .D(n2814), .Y(n3948) );
  OAI21X1 U4972 ( .A(n3949), .B(n2901), .C(n3948), .Y(n4189) );
  XOR2X1 U4973 ( .A(n3950), .B(n4189), .Y(n3951) );
  XNOR2X1 U4974 ( .A(n3952), .B(n3951), .Y(n3957) );
  NAND2X1 U4975 ( .A(n4260), .B(n4189), .Y(n3954) );
  OAI21X1 U4976 ( .A(n4190), .B(n3954), .C(n4045), .Y(n3955) );
  OAI21X1 U4977 ( .A(n4189), .B(n4162), .C(n3955), .Y(n3956) );
  OAI21X1 U4978 ( .A(n4050), .B(n3957), .C(n3956), .Y(inst_EX2MEM_reg_N70) );
  FAX1 U4979 ( .A(n3963), .B(n3959), .C(n3958), .YC(n3939), .YS(n3960) );
  NAND2X1 U4980 ( .A(n4260), .B(n4176), .Y(n3961) );
  OAI21X1 U4981 ( .A(n4177), .B(n3961), .C(n4045), .Y(n3962) );
  OAI21X1 U4982 ( .A(n3963), .B(n4176), .C(n3962), .Y(n3964) );
  OAI21X1 U4983 ( .A(n4050), .B(n3965), .C(n3964), .Y(inst_EX2MEM_reg_N68) );
  FAX1 U4984 ( .A(n4207), .B(n3967), .C(n3966), .YC(n3958), .YS(n3968) );
  NAND2X1 U4985 ( .A(n4150), .B(n4207), .Y(n3969) );
  OAI21X1 U4986 ( .A(n4047), .B(n3969), .C(n4045), .Y(n3970) );
  OAI21X1 U4987 ( .A(n4207), .B(n4150), .C(n3970), .Y(n3971) );
  OAI21X1 U4988 ( .A(n4050), .B(n3972), .C(n3971), .Y(inst_EX2MEM_reg_N67) );
  FAX1 U4989 ( .A(n4151), .B(n3974), .C(n3973), .YC(n3966), .YS(n3975) );
  NAND2X1 U4990 ( .A(n4260), .B(n4171), .Y(n3976) );
  OAI21X1 U4991 ( .A(n4172), .B(n3976), .C(n4045), .Y(n3977) );
  OAI21X1 U4992 ( .A(n4151), .B(n4171), .C(n3977), .Y(n3978) );
  OAI21X1 U4993 ( .A(n4050), .B(n3979), .C(n3978), .Y(inst_EX2MEM_reg_N66) );
  FAX1 U4994 ( .A(n3985), .B(n3981), .C(n3980), .YC(n3973), .YS(n3982) );
  NAND2X1 U4995 ( .A(n4260), .B(n4173), .Y(n3983) );
  OAI21X1 U4996 ( .A(n4174), .B(n3983), .C(n4045), .Y(n3984) );
  OAI21X1 U4997 ( .A(n3985), .B(n4173), .C(n3984), .Y(n3986) );
  OAI21X1 U4998 ( .A(n4033), .B(n3987), .C(n3986), .Y(inst_EX2MEM_reg_N65) );
  FAX1 U4999 ( .A(n3993), .B(n3989), .C(n3988), .YC(n3737), .YS(n3990) );
  NAND2X1 U5000 ( .A(n4260), .B(n4165), .Y(n3991) );
  OAI21X1 U5001 ( .A(n4166), .B(n3991), .C(n4045), .Y(n3992) );
  OAI21X1 U5002 ( .A(n3993), .B(n4165), .C(n3992), .Y(n3994) );
  OAI21X1 U5003 ( .A(n4033), .B(n3995), .C(n3994), .Y(inst_EX2MEM_reg_N63) );
  FAX1 U5004 ( .A(n4060), .B(n3997), .C(n3996), .YC(n3688), .YS(n3998) );
  NAND2X1 U5005 ( .A(n4260), .B(n4060), .Y(n3999) );
  OAI21X1 U5006 ( .A(n4059), .B(n3999), .C(n4045), .Y(n4000) );
  OAI21X1 U5007 ( .A(n4060), .B(n4001), .C(n4000), .Y(n4002) );
  OAI21X1 U5008 ( .A(n4050), .B(n4003), .C(n4002), .Y(inst_EX2MEM_reg_N59) );
  FAX1 U5009 ( .A(n4138), .B(n4005), .C(n4004), .YC(n3677), .YS(n4006) );
  NAND2X1 U5010 ( .A(n4260), .B(n4138), .Y(n4007) );
  OAI21X1 U5011 ( .A(n4139), .B(n4007), .C(n4045), .Y(n4008) );
  OAI21X1 U5012 ( .A(n4138), .B(n4056), .C(n4008), .Y(n4009) );
  OAI21X1 U5013 ( .A(n4050), .B(n4010), .C(n4009), .Y(inst_EX2MEM_reg_N57) );
  FAX1 U5014 ( .A(n4063), .B(n4012), .C(n4011), .YC(n4004), .YS(n4013) );
  NAND2X1 U5015 ( .A(n4260), .B(n4135), .Y(n4014) );
  OAI21X1 U5016 ( .A(n4136), .B(n4014), .C(n4045), .Y(n4015) );
  OAI21X1 U5017 ( .A(n4063), .B(n4135), .C(n4015), .Y(n4016) );
  OAI21X1 U5018 ( .A(n4050), .B(n4017), .C(n4016), .Y(inst_EX2MEM_reg_N56) );
  FAX1 U5019 ( .A(n4023), .B(n4019), .C(n4018), .YC(n2993), .YS(n4020) );
  NAND2X1 U5020 ( .A(n4260), .B(n4104), .Y(n4021) );
  OAI21X1 U5021 ( .A(n4105), .B(n4021), .C(n4045), .Y(n4022) );
  OAI21X1 U5022 ( .A(n4104), .B(n4023), .C(n4022), .Y(n4024) );
  OAI21X1 U5023 ( .A(n4033), .B(n4025), .C(n4024), .Y(inst_EX2MEM_reg_N50) );
  FAX1 U5024 ( .A(n4081), .B(n4027), .C(n4026), .YC(n3571), .YS(n4028) );
  NAND2X1 U5025 ( .A(n4087), .B(n4081), .Y(n4029) );
  OAI21X1 U5026 ( .A(n4047), .B(n4029), .C(n4045), .Y(n4030) );
  OAI21X1 U5027 ( .A(n4087), .B(n4081), .C(n4030), .Y(n4031) );
  OAI21X1 U5028 ( .A(n4033), .B(n4032), .C(n4031), .Y(inst_EX2MEM_reg_N44) );
  FAX1 U5029 ( .A(n4039), .B(n4035), .C(n4034), .YC(n3198), .YS(n4036) );
  INVX1 U5030 ( .A(n4039), .Y(n4076) );
  NAND2X1 U5031 ( .A(n4260), .B(n4075), .Y(n4037) );
  OAI21X1 U5032 ( .A(n4076), .B(n4037), .C(n4045), .Y(n4038) );
  OAI21X1 U5033 ( .A(n4075), .B(n4039), .C(n4038), .Y(n4040) );
  OAI21X1 U5034 ( .A(n4041), .B(n4050), .C(n4040), .Y(inst_EX2MEM_reg_N41) );
  FAX1 U5035 ( .A(n4201), .B(n4043), .C(n4042), .YC(n4034), .YS(n4044) );
  NAND2X1 U5036 ( .A(n4191), .B(n4201), .Y(n4046) );
  OAI21X1 U5037 ( .A(n4047), .B(n4046), .C(n4045), .Y(n4048) );
  OAI21X1 U5038 ( .A(n4191), .B(n4201), .C(n4048), .Y(n4049) );
  OAI21X1 U5039 ( .A(n4051), .B(n4050), .C(n4049), .Y(inst_EX2MEM_reg_N40) );
  NOR2X1 U5040 ( .A(n4258), .B(n4186), .Y(n4255) );
  INVX1 U5041 ( .A(n4160), .Y(n4053) );
  INVX1 U5042 ( .A(n4146), .Y(n4052) );
  AOI22X1 U5043 ( .A(n4053), .B(n4157), .C(n4052), .D(n4143), .Y(n4228) );
  INVX1 U5044 ( .A(n4054), .Y(n4145) );
  OAI22X1 U5045 ( .A(n4059), .B(n4060), .C(n4145), .D(n4144), .Y(n4226) );
  INVX1 U5046 ( .A(n4138), .Y(n4057) );
  INVX1 U5047 ( .A(n4062), .Y(n4055) );
  AOI22X1 U5048 ( .A(n4057), .B(n4056), .C(n4055), .D(n4058), .Y(n4234) );
  AOI22X1 U5049 ( .A(n4062), .B(n4061), .C(n4060), .D(n4059), .Y(n4134) );
  INVX1 U5050 ( .A(n4134), .Y(n4142) );
  INVX1 U5051 ( .A(n4135), .Y(n4064) );
  NOR2X1 U5052 ( .A(n4064), .B(n4063), .Y(n4194) );
  INVX1 U5053 ( .A(n4065), .Y(n4121) );
  AOI22X1 U5054 ( .A(n4121), .B(n4120), .C(n4066), .D(n4124), .Y(n4113) );
  OAI21X1 U5055 ( .A(n4105), .B(n4104), .C(n4113), .Y(n4067) );
  AOI21X1 U5056 ( .A(n4068), .B(n4112), .C(n4067), .Y(n4188) );
  INVX1 U5057 ( .A(n4098), .Y(n4070) );
  INVX1 U5058 ( .A(n4090), .Y(n4069) );
  AOI22X1 U5059 ( .A(n4070), .B(n4095), .C(n4069), .D(n4089), .Y(n4211) );
  INVX1 U5060 ( .A(n4071), .Y(n4082) );
  INVX1 U5061 ( .A(n4072), .Y(n4078) );
  OAI22X1 U5062 ( .A(n4083), .B(n4082), .C(n4077), .D(n4078), .Y(n4214) );
  INVX1 U5063 ( .A(n4258), .Y(n4073) );
  INVX1 U5064 ( .A(n4201), .Y(n4074) );
  AOI22X1 U5065 ( .A(n4073), .B(n4186), .C(n4074), .D(n4191), .Y(n4079) );
  OAI22X1 U5066 ( .A(n4074), .B(n4191), .C(n4076), .D(n4075), .Y(n4239) );
  AOI22X1 U5067 ( .A(n4078), .B(n4077), .C(n4076), .D(n4075), .Y(n4241) );
  OAI21X1 U5068 ( .A(n4079), .B(n4239), .C(n4241), .Y(n4080) );
  INVX1 U5069 ( .A(n4081), .Y(n4088) );
  AOI22X1 U5070 ( .A(n4083), .B(n4082), .C(n4087), .D(n4088), .Y(n4210) );
  OAI21X1 U5071 ( .A(n4214), .B(n4084), .C(n4210), .Y(n4085) );
  INVX1 U5072 ( .A(n4086), .Y(n4093) );
  OAI22X1 U5073 ( .A(n4088), .B(n4087), .C(n4093), .D(n4092), .Y(n4220) );
  INVX1 U5074 ( .A(n4089), .Y(n4091) );
  AOI22X1 U5075 ( .A(n4093), .B(n4092), .C(n4091), .D(n4090), .Y(n4216) );
  OAI21X1 U5076 ( .A(n4094), .B(n4220), .C(n4216), .Y(n4100) );
  INVX1 U5077 ( .A(n4095), .Y(n4097) );
  INVX1 U5078 ( .A(n4096), .Y(n4103) );
  AOI22X1 U5079 ( .A(n4098), .B(n4097), .C(n4102), .D(n4103), .Y(n4212) );
  AOI21X1 U5080 ( .A(n4211), .B(n4100), .C(n4099), .Y(n4108) );
  INVX1 U5081 ( .A(n4101), .Y(n4107) );
  OAI22X1 U5082 ( .A(n4107), .B(n4106), .C(n4103), .D(n4102), .Y(n4215) );
  AOI22X1 U5083 ( .A(n4107), .B(n4106), .C(n4105), .D(n4104), .Y(n4218) );
  OAI21X1 U5084 ( .A(n4108), .B(n4215), .C(n4218), .Y(n4109) );
  NAND2X1 U5085 ( .A(n4188), .B(n4109), .Y(n4133) );
  INVX1 U5086 ( .A(n4110), .Y(n4116) );
  INVX1 U5087 ( .A(n4117), .Y(n4111) );
  NAND2X1 U5088 ( .A(n4111), .B(n4114), .Y(n4122) );
  OAI21X1 U5089 ( .A(n4116), .B(n4115), .C(n4122), .Y(n4238) );
  INVX1 U5090 ( .A(n4112), .Y(n4131) );
  INVX1 U5091 ( .A(n4113), .Y(n4128) );
  NOR2X1 U5092 ( .A(n4121), .B(n4120), .Y(n4123) );
  INVX1 U5093 ( .A(n4114), .Y(n4118) );
  AOI22X1 U5094 ( .A(n4118), .B(n4117), .C(n4116), .D(n4115), .Y(n4119) );
  OAI21X1 U5095 ( .A(n4121), .B(n4120), .C(n4119), .Y(n4244) );
  OAI21X1 U5096 ( .A(n4123), .B(n4122), .C(n4244), .Y(n4127) );
  INVX1 U5097 ( .A(n4124), .Y(n4126) );
  AOI22X1 U5098 ( .A(n4126), .B(n4125), .C(n4131), .D(n4130), .Y(n4236) );
  OAI21X1 U5099 ( .A(n4128), .B(n4127), .C(n4236), .Y(n4129) );
  OAI21X1 U5100 ( .A(n4131), .B(n4130), .C(n4129), .Y(n4132) );
  OAI21X1 U5101 ( .A(n4133), .B(n4238), .C(n4132), .Y(n4140) );
  OAI21X1 U5102 ( .A(n4136), .B(n4135), .C(n4134), .Y(n4137) );
  AOI21X1 U5103 ( .A(n4139), .B(n4138), .C(n4137), .Y(n4245) );
  OAI21X1 U5104 ( .A(n4194), .B(n4140), .C(n4245), .Y(n4141) );
  OAI21X1 U5105 ( .A(n4234), .B(n4142), .C(n4141), .Y(n4148) );
  INVX1 U5106 ( .A(n4143), .Y(n4147) );
  AOI22X1 U5107 ( .A(n4147), .B(n4146), .C(n4145), .D(n4144), .Y(n4227) );
  OAI21X1 U5108 ( .A(n4226), .B(n4148), .C(n4227), .Y(n4156) );
  INVX1 U5109 ( .A(n4149), .Y(n4197) );
  AOI22X1 U5110 ( .A(n4206), .B(n4207), .C(n4152), .D(n4151), .Y(n4153) );
  OAI21X1 U5111 ( .A(n4177), .B(n4176), .C(n4153), .Y(n4179) );
  INVX1 U5112 ( .A(n4179), .Y(n4154) );
  OAI21X1 U5113 ( .A(n4173), .B(n4174), .C(n4154), .Y(n4225) );
  OAI21X1 U5114 ( .A(n4197), .B(n4196), .C(n4155), .Y(n4170) );
  AOI21X1 U5115 ( .A(n4228), .B(n4156), .C(n4170), .Y(n4164) );
  INVX1 U5116 ( .A(n4157), .Y(n4161) );
  AOI22X1 U5117 ( .A(n4190), .B(n4189), .C(n4158), .D(n4167), .Y(n4180) );
  OAI21X1 U5118 ( .A(n4166), .B(n4165), .C(n4180), .Y(n4159) );
  AOI21X1 U5119 ( .A(n4161), .B(n4160), .C(n4159), .Y(n4240) );
  AOI22X1 U5120 ( .A(n4164), .B(n4240), .C(n4163), .D(n4162), .Y(n4185) );
  AOI22X1 U5121 ( .A(n4197), .B(n4196), .C(n4166), .D(n4165), .Y(n4187) );
  INVX1 U5122 ( .A(n4167), .Y(n4169) );
  AOI22X1 U5123 ( .A(n4169), .B(n4168), .C(n4177), .D(n4176), .Y(n4229) );
  OAI21X1 U5124 ( .A(n4187), .B(n4170), .C(n4229), .Y(n4182) );
  AOI22X1 U5125 ( .A(n4174), .B(n4173), .C(n4172), .D(n4171), .Y(n4230) );
  NOR2X1 U5126 ( .A(n4206), .B(n4207), .Y(n4175) );
  OAI21X1 U5127 ( .A(n4177), .B(n4176), .C(n4175), .Y(n4178) );
  OAI21X1 U5128 ( .A(n4230), .B(n4179), .C(n4178), .Y(n4181) );
  OAI21X1 U5129 ( .A(n4182), .B(n4181), .C(n4180), .Y(n4184) );
  AOI21X1 U5130 ( .A(n4185), .B(n4184), .C(n4183), .Y(n4252) );
  AND2X2 U5131 ( .A(n4258), .B(n4186), .Y(n4261) );
  OAI21X1 U5132 ( .A(n4255), .B(n4261), .C(n4187), .Y(n4209) );
  OAI21X1 U5133 ( .A(n4190), .B(n4189), .C(n4188), .Y(n4204) );
  INVX1 U5134 ( .A(n4191), .Y(n4202) );
  NAND3X1 U5135 ( .A(inst_EX2MEM_reg_N6), .B(n4193), .C(n4192), .Y(n4199) );
  OAI21X1 U5136 ( .A(n4197), .B(n4196), .C(n4195), .Y(n4198) );
  NOR2X1 U5137 ( .A(n4199), .B(n4198), .Y(n4200) );
  OAI21X1 U5138 ( .A(n4202), .B(n4201), .C(n4200), .Y(n4203) );
  NOR2X1 U5139 ( .A(n4204), .B(n4203), .Y(n4205) );
  OAI21X1 U5140 ( .A(n4207), .B(n4206), .C(n4205), .Y(n4208) );
  NOR2X1 U5141 ( .A(n4209), .B(n4208), .Y(n4223) );
  NAND3X1 U5142 ( .A(n4212), .B(n4211), .C(n4210), .Y(n4213) );
  NOR2X1 U5143 ( .A(n4214), .B(n4213), .Y(n4222) );
  NAND3X1 U5144 ( .A(n4218), .B(n4217), .C(n4216), .Y(n4219) );
  NOR2X1 U5145 ( .A(n4220), .B(n4219), .Y(n4221) );
  NAND3X1 U5146 ( .A(n4223), .B(n4222), .C(n4221), .Y(n4224) );
  NOR2X1 U5147 ( .A(n4225), .B(n4224), .Y(n4251) );
  INVX1 U5148 ( .A(n4227), .Y(n4232) );
  NAND3X1 U5149 ( .A(n4230), .B(n4229), .C(n4228), .Y(n4231) );
  NOR2X1 U5150 ( .A(n4232), .B(n4231), .Y(n4233) );
  NAND3X1 U5151 ( .A(n4235), .B(n4234), .C(n4233), .Y(n4249) );
  NOR2X1 U5152 ( .A(n4238), .B(n4237), .Y(n4247) );
  NAND3X1 U5153 ( .A(n4242), .B(n4241), .C(n4240), .Y(n4243) );
  NOR2X1 U5154 ( .A(n4244), .B(n4243), .Y(n4246) );
  NAND3X1 U5155 ( .A(n4247), .B(n4246), .C(n4245), .Y(n4248) );
  NOR2X1 U5156 ( .A(n4249), .B(n4248), .Y(n4250) );
  AOI22X1 U5157 ( .A(inst_EX2MEM_reg_N3), .B(n4252), .C(n4251), .D(n4250), .Y(
        n4253) );
  OAI21X1 U5158 ( .A(n4255), .B(n4254), .C(n4253), .Y(n4256) );
  FAX1 U5159 ( .A(n4259), .B(n4258), .C(n4257), .YC(n4042), .YS(n4262) );
  AOI22X1 U5160 ( .A(n4263), .B(n4262), .C(n4261), .D(n4260), .Y(n4264) );
  OAI21X1 U5161 ( .A(op_type_EX[1]), .B(n4265), .C(n4264), .Y(
        inst_EX2MEM_reg_N39) );
  NOR2X1 U5162 ( .A(n2795), .B(n4617), .Y(n4268) );
  AOI22X1 U5163 ( .A(n4294), .B(shifted_address_MEM[0]), .C(n5497), .D(
        jump_inst_addr_MEM[0]), .Y(n4266) );
  OAI21X1 U5164 ( .A(n4268), .B(n4747), .C(n4266), .Y(n2214) );
  AOI22X1 U5165 ( .A(n4294), .B(shifted_address_MEM[1]), .C(n5497), .D(
        jump_inst_addr_MEM[1]), .Y(n4267) );
  OAI21X1 U5166 ( .A(n4268), .B(n4745), .C(n4267), .Y(n2213) );
  OAI21X1 U5167 ( .A(n4312), .B(n5502), .C(n4742), .Y(n4269) );
  AOI22X1 U5168 ( .A(n5497), .B(jump_inst_addr_MEM[3]), .C(n4270), .D(n4269), 
        .Y(n4271) );
  OAI21X1 U5169 ( .A(n4305), .B(n4272), .C(n4271), .Y(n2211) );
  BUFX2 U5170 ( .A(n4727), .Y(n5501) );
  INVX1 U5171 ( .A(n4273), .Y(n4274) );
  OAI21X1 U5172 ( .A(n4274), .B(inst_address[5]), .C(n2795), .Y(n4276) );
  NAND2X1 U5173 ( .A(n5497), .B(jump_inst_addr_MEM[5]), .Y(n4275) );
  OAI21X1 U5174 ( .A(n4280), .B(n4276), .C(n4275), .Y(n4277) );
  AOI21X1 U5175 ( .A(n5526), .B(shifted_address_MEM[5]), .C(n4277), .Y(n4278)
         );
  OAI21X1 U5176 ( .A(n4738), .B(n5501), .C(n4278), .Y(n2209) );
  OAI21X1 U5177 ( .A(n4280), .B(inst_address[6]), .C(n4279), .Y(n4282) );
  NAND2X1 U5178 ( .A(n4294), .B(shifted_address_MEM[6]), .Y(n4281) );
  OAI21X1 U5179 ( .A(n4312), .B(n4282), .C(n4281), .Y(n4283) );
  AOI21X1 U5180 ( .A(n5497), .B(jump_inst_addr_MEM[6]), .C(n4283), .Y(n4284)
         );
  OAI21X1 U5181 ( .A(n4736), .B(n4727), .C(n4284), .Y(n2208) );
  INVX1 U5182 ( .A(inst_address[12]), .Y(n4723) );
  NAND2X1 U5183 ( .A(n5497), .B(jump_inst_addr_MEM[12]), .Y(n4285) );
  OAI21X1 U5184 ( .A(inst_address[12]), .B(n4286), .C(n4285), .Y(n4287) );
  AOI21X1 U5185 ( .A(n5526), .B(shifted_address_MEM[12]), .C(n4287), .Y(n4288)
         );
  OAI21X1 U5186 ( .A(n4289), .B(n4723), .C(n4288), .Y(n2202) );
  AOI21X1 U5187 ( .A(inst_address[12]), .B(n4290), .C(inst_address[13]), .Y(
        n4292) );
  AOI22X1 U5188 ( .A(n4294), .B(shifted_address_MEM[13]), .C(n5497), .D(
        jump_inst_addr_MEM[13]), .Y(n4291) );
  OAI21X1 U5189 ( .A(n4293), .B(n4292), .C(n4291), .Y(n2201) );
  INVX1 U5190 ( .A(inst_address[15]), .Y(n4717) );
  NAND2X1 U5191 ( .A(n4294), .B(shifted_address_MEM[15]), .Y(n4295) );
  OAI21X1 U5192 ( .A(n4296), .B(n4717), .C(n4295), .Y(n4297) );
  AOI21X1 U5193 ( .A(n5497), .B(jump_inst_addr_MEM[15]), .C(n4297), .Y(n4298)
         );
  OAI21X1 U5194 ( .A(inst_address[15]), .B(n4299), .C(n4298), .Y(n2199) );
  OAI21X1 U5195 ( .A(n4301), .B(n4713), .C(n4300), .Y(n4302) );
  AOI21X1 U5196 ( .A(n5497), .B(jump_inst_addr_MEM[17]), .C(n4302), .Y(n4303)
         );
  OAI21X1 U5197 ( .A(n4305), .B(n4304), .C(n4303), .Y(n2197) );
  NOR2X1 U5198 ( .A(instruction_ID[28]), .B(instruction_ID[4]), .Y(n4308) );
  NOR2X1 U5199 ( .A(instruction_ID[26]), .B(instruction_ID[31]), .Y(n4309) );
  NOR2X1 U5200 ( .A(instruction_ID[27]), .B(instruction_ID[30]), .Y(n4306) );
  NAND2X1 U5201 ( .A(n4309), .B(n4306), .Y(n4330) );
  NOR2X1 U5202 ( .A(instruction_ID[29]), .B(n4330), .Y(n4307) );
  NAND3X1 U5203 ( .A(inst_ID2EX_reg_N108), .B(n4308), .C(n4307), .Y(n4324) );
  NOR2X1 U5204 ( .A(instruction_ID[0]), .B(n4324), .Y(n4314) );
  NAND2X1 U5205 ( .A(n4314), .B(n4676), .Y(n4318) );
  INVX1 U5206 ( .A(instruction_ID[28]), .Y(n4626) );
  INVX1 U5207 ( .A(instruction_ID[30]), .Y(n4622) );
  NAND3X1 U5208 ( .A(instruction_ID[27]), .B(n4626), .C(n4622), .Y(n4311) );
  NOR2X1 U5209 ( .A(instruction_ID[29]), .B(n5524), .Y(n4326) );
  NAND2X1 U5210 ( .A(n4326), .B(n4309), .Y(n4310) );
  NOR2X1 U5211 ( .A(n4311), .B(n4310), .Y(n4327) );
  INVX1 U5212 ( .A(instruction_ID[29]), .Y(n4624) );
  NOR2X1 U5213 ( .A(n4312), .B(n4311), .Y(n4313) );
  NAND3X1 U5214 ( .A(instruction_ID[26]), .B(instruction_ID[31]), .C(n4313), 
        .Y(n4321) );
  NOR2X1 U5215 ( .A(instruction_ID[2]), .B(n4680), .Y(n4317) );
  NAND3X1 U5216 ( .A(instruction_ID[3]), .B(n4314), .C(n4317), .Y(n4322) );
  OAI21X1 U5217 ( .A(n4624), .B(n4321), .C(n4322), .Y(n4315) );
  NOR2X1 U5218 ( .A(n4327), .B(n4315), .Y(n4316) );
  OAI21X1 U5219 ( .A(instruction_ID[1]), .B(n4318), .C(n4316), .Y(
        inst_ID2EX_reg_N3) );
  AOI21X1 U5220 ( .A(instruction_ID[2]), .B(n4680), .C(n4317), .Y(n4319) );
  OAI21X1 U5221 ( .A(n4319), .B(n4318), .C(n4321), .Y(inst_ID2EX_reg_N4) );
  NOR2X1 U5222 ( .A(instruction_ID[1]), .B(n4678), .Y(n4320) );
  NAND3X1 U5223 ( .A(instruction_ID[0]), .B(n4320), .C(n4676), .Y(n4325) );
  AND2X2 U5224 ( .A(n4322), .B(n4321), .Y(n4323) );
  OAI21X1 U5225 ( .A(n4325), .B(n4324), .C(n4323), .Y(inst_ID2EX_reg_N5) );
  NAND2X1 U5226 ( .A(n4326), .B(instruction_ID[28]), .Y(n4329) );
  OAI21X1 U5227 ( .A(n4330), .B(n4329), .C(n4328), .Y(inst_ID2EX_reg_N6) );
  OAI21X1 U5228 ( .A(inst_addr_EX[2]), .B(n4332), .C(n4426), .Y(n4331) );
  AOI21X1 U5229 ( .A(inst_addr_EX[2]), .B(n4332), .C(n4331), .Y(
        inst_EX2MEM_reg_N9) );
  INVX1 U5230 ( .A(n4333), .Y(n4334) );
  NOR2X1 U5231 ( .A(n4335), .B(n4334), .Y(n4337) );
  OAI21X1 U5232 ( .A(inst_addr_EX[3]), .B(n4337), .C(n4426), .Y(n4336) );
  AOI21X1 U5233 ( .A(inst_addr_EX[3]), .B(n4337), .C(n4336), .Y(
        inst_EX2MEM_reg_N10) );
  INVX1 U5234 ( .A(n4338), .Y(n4339) );
  NOR2X1 U5235 ( .A(n4340), .B(n4339), .Y(n4342) );
  OAI21X1 U5236 ( .A(inst_addr_EX[4]), .B(n4342), .C(n4426), .Y(n4341) );
  AOI21X1 U5237 ( .A(inst_addr_EX[4]), .B(n4342), .C(n4341), .Y(
        inst_EX2MEM_reg_N11) );
  INVX1 U5238 ( .A(n4343), .Y(n4344) );
  NOR2X1 U5239 ( .A(n4345), .B(n4344), .Y(n4347) );
  OAI21X1 U5240 ( .A(inst_addr_EX[5]), .B(n4347), .C(n4426), .Y(n4346) );
  AOI21X1 U5241 ( .A(inst_addr_EX[5]), .B(n4347), .C(n4346), .Y(
        inst_EX2MEM_reg_N12) );
  INVX1 U5242 ( .A(n4348), .Y(n4349) );
  NOR2X1 U5243 ( .A(n4350), .B(n4349), .Y(n4352) );
  OAI21X1 U5244 ( .A(inst_addr_EX[6]), .B(n4352), .C(n4426), .Y(n4351) );
  AOI21X1 U5245 ( .A(inst_addr_EX[6]), .B(n4352), .C(n4351), .Y(
        inst_EX2MEM_reg_N13) );
  INVX1 U5246 ( .A(n4353), .Y(n4354) );
  NOR2X1 U5247 ( .A(n4355), .B(n4354), .Y(n4357) );
  OAI21X1 U5248 ( .A(inst_addr_EX[7]), .B(n4357), .C(n4426), .Y(n4356) );
  AOI21X1 U5249 ( .A(inst_addr_EX[7]), .B(n4357), .C(n4356), .Y(
        inst_EX2MEM_reg_N14) );
  NOR2X1 U5250 ( .A(n4359), .B(n4358), .Y(n4361) );
  OAI21X1 U5251 ( .A(inst_addr_EX[8]), .B(n4361), .C(n4426), .Y(n4360) );
  AOI21X1 U5252 ( .A(inst_addr_EX[8]), .B(n4361), .C(n4360), .Y(
        inst_EX2MEM_reg_N15) );
  AOI21X1 U5253 ( .A(n4363), .B(jump_inst_addr_EX[8]), .C(n4362), .Y(n4365) );
  OAI21X1 U5254 ( .A(inst_addr_EX[10]), .B(n4365), .C(n4426), .Y(n4364) );
  AOI21X1 U5255 ( .A(inst_addr_EX[10]), .B(n4365), .C(n4364), .Y(
        inst_EX2MEM_reg_N17) );
  MUX2X1 U5256 ( .B(n4367), .A(jump_inst_addr_EX[9]), .S(n4366), .Y(n4369) );
  OAI21X1 U5257 ( .A(inst_addr_EX[11]), .B(n4369), .C(n4426), .Y(n4368) );
  AOI21X1 U5258 ( .A(inst_addr_EX[11]), .B(n4369), .C(n4368), .Y(
        inst_EX2MEM_reg_N18) );
  AOI21X1 U5259 ( .A(n4371), .B(jump_inst_addr_EX[11]), .C(n4370), .Y(n4373)
         );
  OAI21X1 U5260 ( .A(inst_addr_EX[13]), .B(n4373), .C(n4426), .Y(n4372) );
  AOI21X1 U5261 ( .A(inst_addr_EX[13]), .B(n4373), .C(n4372), .Y(
        inst_EX2MEM_reg_N20) );
  MUX2X1 U5262 ( .B(n4375), .A(jump_inst_addr_EX[12]), .S(n4374), .Y(n4377) );
  OAI21X1 U5263 ( .A(inst_addr_EX[14]), .B(n4377), .C(n4426), .Y(n4376) );
  AOI21X1 U5264 ( .A(inst_addr_EX[14]), .B(n4377), .C(n4376), .Y(
        inst_EX2MEM_reg_N21) );
  AOI21X1 U5265 ( .A(n4379), .B(jump_inst_addr_EX[14]), .C(n4378), .Y(n4381)
         );
  OAI21X1 U5266 ( .A(inst_addr_EX[16]), .B(n4381), .C(n4426), .Y(n4380) );
  AOI21X1 U5267 ( .A(inst_addr_EX[16]), .B(n4381), .C(n4380), .Y(
        inst_EX2MEM_reg_N23) );
  MUX2X1 U5268 ( .B(n4419), .A(n4414), .S(n4382), .Y(n4384) );
  OAI21X1 U5269 ( .A(inst_addr_EX[17]), .B(n4384), .C(n4426), .Y(n4383) );
  AOI21X1 U5270 ( .A(inst_addr_EX[17]), .B(n4384), .C(n4383), .Y(
        inst_EX2MEM_reg_N24) );
  AOI21X1 U5271 ( .A(n4386), .B(n4414), .C(n4385), .Y(n4388) );
  OAI21X1 U5272 ( .A(inst_addr_EX[19]), .B(n4388), .C(n4426), .Y(n4387) );
  AOI21X1 U5273 ( .A(inst_addr_EX[19]), .B(n4388), .C(n4387), .Y(
        inst_EX2MEM_reg_N26) );
  OAI21X1 U5274 ( .A(n4414), .B(n4390), .C(n4389), .Y(n4392) );
  OAI21X1 U5275 ( .A(n4393), .B(n4392), .C(n4426), .Y(n4391) );
  AOI21X1 U5276 ( .A(n4393), .B(n4392), .C(n4391), .Y(inst_EX2MEM_reg_N28) );
  AOI21X1 U5277 ( .A(n4414), .B(n4395), .C(n4394), .Y(n4397) );
  OAI21X1 U5278 ( .A(inst_addr_EX[22]), .B(n4397), .C(n4426), .Y(n4396) );
  AOI21X1 U5279 ( .A(inst_addr_EX[22]), .B(n4397), .C(n4396), .Y(
        inst_EX2MEM_reg_N29) );
  AND2X2 U5280 ( .A(n4399), .B(n4398), .Y(n4401) );
  OAI21X1 U5281 ( .A(inst_addr_EX[23]), .B(n4401), .C(n4426), .Y(n4400) );
  AOI21X1 U5282 ( .A(inst_addr_EX[23]), .B(n4401), .C(n4400), .Y(
        inst_EX2MEM_reg_N30) );
  OAI21X1 U5283 ( .A(n4414), .B(n4403), .C(n4402), .Y(n4405) );
  OAI21X1 U5284 ( .A(n4406), .B(n4405), .C(n4426), .Y(n4404) );
  AOI21X1 U5285 ( .A(n4406), .B(n4405), .C(n4404), .Y(inst_EX2MEM_reg_N33) );
  NOR2X1 U5286 ( .A(n4408), .B(n4407), .Y(n4410) );
  OAI21X1 U5287 ( .A(inst_addr_EX[27]), .B(n4410), .C(n4426), .Y(n4409) );
  AOI21X1 U5288 ( .A(inst_addr_EX[27]), .B(n4410), .C(n4409), .Y(
        inst_EX2MEM_reg_N34) );
  FAX1 U5289 ( .A(inst_addr_EX[28]), .B(n4414), .C(n4411), .YC(n4425), .YS(
        n3650) );
  NAND2X1 U5290 ( .A(n4414), .B(n4425), .Y(n4415) );
  OAI21X1 U5291 ( .A(n4414), .B(n4425), .C(n4415), .Y(n4413) );
  OAI21X1 U5292 ( .A(n4420), .B(n4413), .C(n4426), .Y(n4412) );
  AOI21X1 U5293 ( .A(n4420), .B(n4413), .C(n4412), .Y(inst_EX2MEM_reg_N36) );
  OAI21X1 U5294 ( .A(n4414), .B(n4425), .C(inst_addr_EX[29]), .Y(n4422) );
  NAND2X1 U5295 ( .A(n4415), .B(n4422), .Y(n4418) );
  NAND2X1 U5296 ( .A(inst_addr_EX[30]), .B(n4419), .Y(n4423) );
  OAI21X1 U5297 ( .A(inst_addr_EX[30]), .B(n4419), .C(n4423), .Y(n4417) );
  OAI21X1 U5298 ( .A(n4418), .B(n4417), .C(n4426), .Y(n4416) );
  AOI21X1 U5299 ( .A(n4418), .B(n4417), .C(n4416), .Y(inst_EX2MEM_reg_N37) );
  NOR2X1 U5300 ( .A(inst_addr_EX[30]), .B(n4419), .Y(n4421) );
  NAND2X1 U5301 ( .A(n4421), .B(n4420), .Y(n4424) );
  OAI22X1 U5302 ( .A(n4425), .B(n4424), .C(n4423), .D(n4422), .Y(n4428) );
  OAI21X1 U5303 ( .A(inst_addr_EX[31]), .B(n4428), .C(n4426), .Y(n4427) );
  AOI21X1 U5304 ( .A(inst_addr_EX[31]), .B(n4428), .C(n4427), .Y(
        inst_EX2MEM_reg_N38) );
  NOR2X1 U5305 ( .A(op_type_MEM[3]), .B(n4429), .Y(n4431) );
  NAND3X1 U5306 ( .A(u_MEM2WB_reg_N4), .B(n4431), .C(n4430), .Y(n4445) );
  NOR2X1 U5307 ( .A(alu_result_MEM[1]), .B(n4432), .Y(n4444) );
  NAND2X1 U5308 ( .A(alu_result_MEM[0]), .B(n4444), .Y(n4885) );
  NOR2X1 U5309 ( .A(n4445), .B(n4885), .Y(n4526) );
  AOI22X1 U5310 ( .A(inst_data_MEM_data[160]), .B(n4526), .C(
        inst_data_MEM_data[224]), .D(n2797), .Y(n4450) );
  NOR2X1 U5311 ( .A(alu_result_MEM[2]), .B(n4434), .Y(n4438) );
  NAND2X1 U5312 ( .A(n4438), .B(n4443), .Y(n4757) );
  NOR2X1 U5313 ( .A(n4445), .B(n4757), .Y(n4602) );
  INVX1 U5314 ( .A(n4795), .Y(n4436) );
  NOR2X1 U5315 ( .A(n4436), .B(n4445), .Y(n4603) );
  AOI22X1 U5316 ( .A(inst_data_MEM_data[64]), .B(n4435), .C(
        inst_data_MEM_data[32]), .D(n4437), .Y(n4449) );
  NAND2X1 U5317 ( .A(alu_result_MEM[0]), .B(n4438), .Y(n4750) );
  NAND2X1 U5318 ( .A(n4439), .B(n4443), .Y(n4875) );
  AOI22X1 U5319 ( .A(inst_data_MEM_data[96]), .B(n2799), .C(
        inst_data_MEM_data[192]), .D(n2800), .Y(n4447) );
  NAND2X1 U5320 ( .A(n4441), .B(n4443), .Y(n4833) );
  NOR2X1 U5321 ( .A(n4833), .B(n4445), .Y(n4609) );
  NAND2X1 U5322 ( .A(n4444), .B(n4443), .Y(n4926) );
  AOI22X1 U5323 ( .A(inst_data_MEM_data[0]), .B(n4442), .C(
        inst_data_MEM_data[128]), .D(n2798), .Y(n4446) );
  AND2X2 U5324 ( .A(n4447), .B(n4446), .Y(n4448) );
  NAND3X1 U5325 ( .A(n4450), .B(n4449), .C(n4448), .Y(u_MEM2WB_reg_N7) );
  AOI22X1 U5326 ( .A(n2798), .B(inst_data_MEM_data[129]), .C(n4451), .D(
        inst_data_MEM_data[161]), .Y(n4456) );
  AOI22X1 U5327 ( .A(n4435), .B(inst_data_MEM_data[65]), .C(n2797), .D(
        inst_data_MEM_data[225]), .Y(n4455) );
  AOI22X1 U5328 ( .A(n2799), .B(inst_data_MEM_data[97]), .C(n4603), .D(
        inst_data_MEM_data[33]), .Y(n4453) );
  AOI22X1 U5329 ( .A(n4442), .B(inst_data_MEM_data[1]), .C(n2800), .D(
        inst_data_MEM_data[193]), .Y(n4452) );
  AND2X2 U5330 ( .A(n4453), .B(n4452), .Y(n4454) );
  NAND3X1 U5331 ( .A(n4456), .B(n4455), .C(n4454), .Y(u_MEM2WB_reg_N8) );
  AOI22X1 U5332 ( .A(n2799), .B(inst_data_MEM_data[98]), .C(n2797), .D(
        inst_data_MEM_data[226]), .Y(n4462) );
  AOI22X1 U5333 ( .A(n4442), .B(inst_data_MEM_data[2]), .C(n4437), .D(
        inst_data_MEM_data[34]), .Y(n4461) );
  AOI22X1 U5334 ( .A(n4435), .B(inst_data_MEM_data[66]), .C(n4451), .D(
        inst_data_MEM_data[162]), .Y(n4459) );
  AOI22X1 U5335 ( .A(n2798), .B(inst_data_MEM_data[130]), .C(n2800), .D(
        inst_data_MEM_data[194]), .Y(n4458) );
  AND2X2 U5336 ( .A(n4459), .B(n4458), .Y(n4460) );
  NAND3X1 U5337 ( .A(n4462), .B(n4461), .C(n4460), .Y(u_MEM2WB_reg_N9) );
  AOI22X1 U5338 ( .A(n4435), .B(inst_data_MEM_data[67]), .C(n4437), .D(
        inst_data_MEM_data[35]), .Y(n4467) );
  AOI22X1 U5339 ( .A(n4526), .B(inst_data_MEM_data[163]), .C(n2797), .D(
        inst_data_MEM_data[227]), .Y(n4466) );
  AOI22X1 U5340 ( .A(n4442), .B(inst_data_MEM_data[3]), .C(n2799), .D(
        inst_data_MEM_data[99]), .Y(n4464) );
  AOI22X1 U5341 ( .A(n2798), .B(inst_data_MEM_data[131]), .C(n2800), .D(
        inst_data_MEM_data[195]), .Y(n4463) );
  AND2X2 U5342 ( .A(n4464), .B(n4463), .Y(n4465) );
  NAND3X1 U5343 ( .A(n4467), .B(n4466), .C(n4465), .Y(u_MEM2WB_reg_N10) );
  AOI22X1 U5344 ( .A(n2800), .B(inst_data_MEM_data[196]), .C(n4526), .D(
        inst_data_MEM_data[164]), .Y(n4473) );
  AOI22X1 U5345 ( .A(n4435), .B(inst_data_MEM_data[68]), .C(n2797), .D(
        inst_data_MEM_data[228]), .Y(n4472) );
  AOI22X1 U5346 ( .A(n4442), .B(inst_data_MEM_data[4]), .C(n4437), .D(
        inst_data_MEM_data[36]), .Y(n4470) );
  AOI22X1 U5347 ( .A(n2798), .B(inst_data_MEM_data[132]), .C(n2799), .D(
        inst_data_MEM_data[100]), .Y(n4469) );
  AND2X2 U5348 ( .A(n4470), .B(n4469), .Y(n4471) );
  NAND3X1 U5349 ( .A(n4473), .B(n4472), .C(n4471), .Y(u_MEM2WB_reg_N11) );
  AOI22X1 U5350 ( .A(n2799), .B(inst_data_MEM_data[101]), .C(n2797), .D(
        inst_data_MEM_data[229]), .Y(n4479) );
  AOI22X1 U5351 ( .A(n4442), .B(inst_data_MEM_data[5]), .C(n4451), .D(
        inst_data_MEM_data[165]), .Y(n4478) );
  AOI22X1 U5352 ( .A(n4435), .B(inst_data_MEM_data[69]), .C(n4437), .D(
        inst_data_MEM_data[37]), .Y(n4476) );
  AOI22X1 U5353 ( .A(n2798), .B(inst_data_MEM_data[133]), .C(n2800), .D(
        inst_data_MEM_data[197]), .Y(n4475) );
  AND2X2 U5354 ( .A(n4476), .B(n4475), .Y(n4477) );
  NAND3X1 U5355 ( .A(n4479), .B(n4478), .C(n4477), .Y(u_MEM2WB_reg_N12) );
  AOI22X1 U5356 ( .A(n2800), .B(inst_data_MEM_data[198]), .C(n4526), .D(
        inst_data_MEM_data[166]), .Y(n4484) );
  AOI22X1 U5357 ( .A(n2799), .B(inst_data_MEM_data[102]), .C(n4435), .D(
        inst_data_MEM_data[70]), .Y(n4483) );
  AOI22X1 U5358 ( .A(n4442), .B(inst_data_MEM_data[6]), .C(n2798), .D(
        inst_data_MEM_data[134]), .Y(n4481) );
  AOI22X1 U5359 ( .A(n4437), .B(inst_data_MEM_data[38]), .C(n2797), .D(
        inst_data_MEM_data[230]), .Y(n4480) );
  AND2X2 U5360 ( .A(n4481), .B(n4480), .Y(n4482) );
  NAND3X1 U5361 ( .A(n4484), .B(n4483), .C(n4482), .Y(u_MEM2WB_reg_N13) );
  AOI22X1 U5362 ( .A(n4442), .B(inst_data_MEM_data[7]), .C(n4437), .D(
        inst_data_MEM_data[39]), .Y(n4489) );
  AOI22X1 U5363 ( .A(n2799), .B(inst_data_MEM_data[103]), .C(n2800), .D(
        inst_data_MEM_data[199]), .Y(n4488) );
  AOI22X1 U5364 ( .A(n2798), .B(inst_data_MEM_data[135]), .C(n4526), .D(
        inst_data_MEM_data[167]), .Y(n4486) );
  AOI22X1 U5365 ( .A(n4435), .B(inst_data_MEM_data[71]), .C(n2797), .D(
        inst_data_MEM_data[231]), .Y(n4485) );
  AND2X2 U5366 ( .A(n4486), .B(n4485), .Y(n4487) );
  NAND3X1 U5367 ( .A(n4489), .B(n4488), .C(n4487), .Y(u_MEM2WB_reg_N14) );
  AOI22X1 U5368 ( .A(n2799), .B(inst_data_MEM_data[104]), .C(n2797), .D(
        inst_data_MEM_data[232]), .Y(n4494) );
  AOI22X1 U5369 ( .A(n4435), .B(inst_data_MEM_data[72]), .C(n4437), .D(
        inst_data_MEM_data[40]), .Y(n4493) );
  AOI22X1 U5370 ( .A(n2800), .B(inst_data_MEM_data[200]), .C(n4526), .D(
        inst_data_MEM_data[168]), .Y(n4491) );
  AOI22X1 U5371 ( .A(n4442), .B(inst_data_MEM_data[8]), .C(n2798), .D(
        inst_data_MEM_data[136]), .Y(n4490) );
  AND2X2 U5372 ( .A(n4491), .B(n4490), .Y(n4492) );
  NAND3X1 U5373 ( .A(n4494), .B(n4493), .C(n4492), .Y(u_MEM2WB_reg_N15) );
  AOI22X1 U5374 ( .A(n4442), .B(inst_data_MEM_data[9]), .C(n2798), .D(
        inst_data_MEM_data[137]), .Y(n4499) );
  AOI22X1 U5375 ( .A(n2799), .B(inst_data_MEM_data[105]), .C(n2797), .D(
        inst_data_MEM_data[233]), .Y(n4498) );
  AOI22X1 U5376 ( .A(n2800), .B(inst_data_MEM_data[201]), .C(n4435), .D(
        inst_data_MEM_data[73]), .Y(n4496) );
  AOI22X1 U5377 ( .A(n4437), .B(inst_data_MEM_data[41]), .C(n4451), .D(
        inst_data_MEM_data[169]), .Y(n4495) );
  AND2X2 U5378 ( .A(n4496), .B(n4495), .Y(n4497) );
  NAND3X1 U5379 ( .A(n4499), .B(n4498), .C(n4497), .Y(u_MEM2WB_reg_N16) );
  AOI22X1 U5380 ( .A(n4442), .B(inst_data_MEM_data[10]), .C(n2800), .D(
        inst_data_MEM_data[202]), .Y(n4504) );
  AOI22X1 U5381 ( .A(n2798), .B(inst_data_MEM_data[138]), .C(n2797), .D(
        inst_data_MEM_data[234]), .Y(n4503) );
  AOI22X1 U5382 ( .A(n2799), .B(inst_data_MEM_data[106]), .C(n4435), .D(
        inst_data_MEM_data[74]), .Y(n4501) );
  AOI22X1 U5383 ( .A(n4437), .B(inst_data_MEM_data[42]), .C(n4526), .D(
        inst_data_MEM_data[170]), .Y(n4500) );
  AND2X2 U5384 ( .A(n4501), .B(n4500), .Y(n4502) );
  NAND3X1 U5385 ( .A(n4504), .B(n4503), .C(n4502), .Y(u_MEM2WB_reg_N17) );
  AOI22X1 U5386 ( .A(n2798), .B(inst_data_MEM_data[139]), .C(n4435), .D(
        inst_data_MEM_data[75]), .Y(n4509) );
  AOI22X1 U5387 ( .A(n2799), .B(inst_data_MEM_data[107]), .C(n4451), .D(
        inst_data_MEM_data[171]), .Y(n4508) );
  AOI22X1 U5388 ( .A(n4442), .B(inst_data_MEM_data[11]), .C(n2797), .D(
        inst_data_MEM_data[235]), .Y(n4506) );
  AOI22X1 U5389 ( .A(n2800), .B(inst_data_MEM_data[203]), .C(n4437), .D(
        inst_data_MEM_data[43]), .Y(n4505) );
  AND2X2 U5390 ( .A(n4506), .B(n4505), .Y(n4507) );
  NAND3X1 U5391 ( .A(n4509), .B(n4508), .C(n4507), .Y(u_MEM2WB_reg_N18) );
  AOI22X1 U5392 ( .A(n4603), .B(inst_data_MEM_data[44]), .C(n2797), .D(
        inst_data_MEM_data[236]), .Y(n4514) );
  AOI22X1 U5393 ( .A(n2798), .B(inst_data_MEM_data[140]), .C(n2800), .D(
        inst_data_MEM_data[204]), .Y(n4513) );
  AOI22X1 U5394 ( .A(n2799), .B(inst_data_MEM_data[108]), .C(n4526), .D(
        inst_data_MEM_data[172]), .Y(n4511) );
  AOI22X1 U5395 ( .A(n4442), .B(inst_data_MEM_data[12]), .C(n4435), .D(
        inst_data_MEM_data[76]), .Y(n4510) );
  AND2X2 U5396 ( .A(n4511), .B(n4510), .Y(n4512) );
  NAND3X1 U5397 ( .A(n4514), .B(n4513), .C(n4512), .Y(u_MEM2WB_reg_N19) );
  AOI22X1 U5398 ( .A(n4609), .B(inst_data_MEM_data[13]), .C(n2797), .D(
        inst_data_MEM_data[237]), .Y(n4520) );
  AOI22X1 U5399 ( .A(n4435), .B(inst_data_MEM_data[77]), .C(n4451), .D(
        inst_data_MEM_data[173]), .Y(n4519) );
  AOI22X1 U5400 ( .A(n2799), .B(inst_data_MEM_data[109]), .C(n4603), .D(
        inst_data_MEM_data[45]), .Y(n4517) );
  AOI22X1 U5401 ( .A(n2798), .B(inst_data_MEM_data[141]), .C(n2800), .D(
        inst_data_MEM_data[205]), .Y(n4516) );
  AND2X2 U5402 ( .A(n4517), .B(n4516), .Y(n4518) );
  NAND3X1 U5403 ( .A(n4520), .B(n4519), .C(n4518), .Y(u_MEM2WB_reg_N20) );
  AOI22X1 U5404 ( .A(n4437), .B(inst_data_MEM_data[46]), .C(n4526), .D(
        inst_data_MEM_data[174]), .Y(n4525) );
  AOI22X1 U5405 ( .A(n4435), .B(inst_data_MEM_data[78]), .C(n2797), .D(
        inst_data_MEM_data[238]), .Y(n4524) );
  AOI22X1 U5406 ( .A(n4442), .B(inst_data_MEM_data[14]), .C(n2799), .D(
        inst_data_MEM_data[110]), .Y(n4522) );
  AOI22X1 U5407 ( .A(n2798), .B(inst_data_MEM_data[142]), .C(n2800), .D(
        inst_data_MEM_data[206]), .Y(n4521) );
  AND2X2 U5408 ( .A(n4522), .B(n4521), .Y(n4523) );
  NAND3X1 U5409 ( .A(n4525), .B(n4524), .C(n4523), .Y(u_MEM2WB_reg_N21) );
  AOI22X1 U5410 ( .A(n2800), .B(inst_data_MEM_data[207]), .C(n4437), .D(
        inst_data_MEM_data[47]), .Y(n4531) );
  AOI22X1 U5411 ( .A(n2798), .B(inst_data_MEM_data[143]), .C(n4435), .D(
        inst_data_MEM_data[79]), .Y(n4530) );
  AOI22X1 U5412 ( .A(n4609), .B(inst_data_MEM_data[15]), .C(n4526), .D(
        inst_data_MEM_data[175]), .Y(n4528) );
  AOI22X1 U5413 ( .A(n2799), .B(inst_data_MEM_data[111]), .C(n2797), .D(
        inst_data_MEM_data[239]), .Y(n4527) );
  AND2X2 U5414 ( .A(n4528), .B(n4527), .Y(n4529) );
  NAND3X1 U5415 ( .A(n4531), .B(n4530), .C(n4529), .Y(u_MEM2WB_reg_N22) );
  AOI22X1 U5416 ( .A(n4451), .B(inst_data_MEM_data[176]), .C(n2797), .D(
        inst_data_MEM_data[240]), .Y(n4536) );
  AOI22X1 U5417 ( .A(n2798), .B(inst_data_MEM_data[144]), .C(n2800), .D(
        inst_data_MEM_data[208]), .Y(n4535) );
  AOI22X1 U5418 ( .A(n4609), .B(inst_data_MEM_data[16]), .C(n4435), .D(
        inst_data_MEM_data[80]), .Y(n4533) );
  AOI22X1 U5419 ( .A(n2799), .B(inst_data_MEM_data[112]), .C(n4603), .D(
        inst_data_MEM_data[48]), .Y(n4532) );
  AND2X2 U5420 ( .A(n4533), .B(n4532), .Y(n4534) );
  NAND3X1 U5421 ( .A(n4536), .B(n4535), .C(n4534), .Y(u_MEM2WB_reg_N23) );
  AOI22X1 U5422 ( .A(n4609), .B(inst_data_MEM_data[17]), .C(n2800), .D(
        inst_data_MEM_data[209]), .Y(n4541) );
  AOI22X1 U5423 ( .A(n2798), .B(inst_data_MEM_data[145]), .C(n4602), .D(
        inst_data_MEM_data[81]), .Y(n4540) );
  AOI22X1 U5424 ( .A(n2799), .B(inst_data_MEM_data[113]), .C(n2797), .D(
        inst_data_MEM_data[241]), .Y(n4538) );
  AOI22X1 U5425 ( .A(n4437), .B(inst_data_MEM_data[49]), .C(n4451), .D(
        inst_data_MEM_data[177]), .Y(n4537) );
  AND2X2 U5426 ( .A(n4538), .B(n4537), .Y(n4539) );
  NAND3X1 U5427 ( .A(n4541), .B(n4540), .C(n4539), .Y(u_MEM2WB_reg_N24) );
  AOI22X1 U5428 ( .A(n4435), .B(inst_data_MEM_data[82]), .C(n4437), .D(
        inst_data_MEM_data[50]), .Y(n4546) );
  AOI22X1 U5429 ( .A(n2800), .B(inst_data_MEM_data[210]), .C(n2797), .D(
        inst_data_MEM_data[242]), .Y(n4545) );
  AOI22X1 U5430 ( .A(n4609), .B(inst_data_MEM_data[18]), .C(n2798), .D(
        inst_data_MEM_data[146]), .Y(n4543) );
  AOI22X1 U5431 ( .A(n2799), .B(inst_data_MEM_data[114]), .C(n4451), .D(
        inst_data_MEM_data[178]), .Y(n4542) );
  AND2X2 U5432 ( .A(n4543), .B(n4542), .Y(n4544) );
  NAND3X1 U5433 ( .A(n4546), .B(n4545), .C(n4544), .Y(u_MEM2WB_reg_N25) );
  AOI22X1 U5434 ( .A(n2800), .B(inst_data_MEM_data[211]), .C(n4602), .D(
        inst_data_MEM_data[83]), .Y(n4551) );
  AOI22X1 U5435 ( .A(n2798), .B(inst_data_MEM_data[147]), .C(n2799), .D(
        inst_data_MEM_data[115]), .Y(n4550) );
  AOI22X1 U5436 ( .A(n4437), .B(inst_data_MEM_data[51]), .C(n2797), .D(
        inst_data_MEM_data[243]), .Y(n4548) );
  AOI22X1 U5437 ( .A(n4442), .B(inst_data_MEM_data[19]), .C(n4451), .D(
        inst_data_MEM_data[179]), .Y(n4547) );
  AND2X2 U5438 ( .A(n4548), .B(n4547), .Y(n4549) );
  NAND3X1 U5439 ( .A(n4551), .B(n4550), .C(n4549), .Y(u_MEM2WB_reg_N26) );
  AOI22X1 U5440 ( .A(n2799), .B(inst_data_MEM_data[116]), .C(n2797), .D(
        inst_data_MEM_data[244]), .Y(n4556) );
  AOI22X1 U5441 ( .A(n2800), .B(inst_data_MEM_data[212]), .C(n4603), .D(
        inst_data_MEM_data[52]), .Y(n4555) );
  AOI22X1 U5442 ( .A(n4609), .B(inst_data_MEM_data[20]), .C(n4602), .D(
        inst_data_MEM_data[84]), .Y(n4553) );
  AOI22X1 U5443 ( .A(n2798), .B(inst_data_MEM_data[148]), .C(n4451), .D(
        inst_data_MEM_data[180]), .Y(n4552) );
  AND2X2 U5444 ( .A(n4553), .B(n4552), .Y(n4554) );
  NAND3X1 U5445 ( .A(n4556), .B(n4555), .C(n4554), .Y(u_MEM2WB_reg_N27) );
  AOI22X1 U5446 ( .A(n2800), .B(inst_data_MEM_data[213]), .C(n4602), .D(
        inst_data_MEM_data[85]), .Y(n4561) );
  AOI22X1 U5447 ( .A(n2798), .B(inst_data_MEM_data[149]), .C(n4603), .D(
        inst_data_MEM_data[53]), .Y(n4560) );
  AOI22X1 U5448 ( .A(n4609), .B(inst_data_MEM_data[21]), .C(n2797), .D(
        inst_data_MEM_data[245]), .Y(n4558) );
  AOI22X1 U5449 ( .A(n2799), .B(inst_data_MEM_data[117]), .C(n4451), .D(
        inst_data_MEM_data[181]), .Y(n4557) );
  AND2X2 U5450 ( .A(n4558), .B(n4557), .Y(n4559) );
  NAND3X1 U5451 ( .A(n4561), .B(n4560), .C(n4559), .Y(u_MEM2WB_reg_N28) );
  AOI22X1 U5452 ( .A(n2800), .B(inst_data_MEM_data[214]), .C(n4602), .D(
        inst_data_MEM_data[86]), .Y(n4566) );
  AOI22X1 U5453 ( .A(n4442), .B(inst_data_MEM_data[22]), .C(n2798), .D(
        inst_data_MEM_data[150]), .Y(n4565) );
  AOI22X1 U5454 ( .A(n4437), .B(inst_data_MEM_data[54]), .C(n2797), .D(
        inst_data_MEM_data[246]), .Y(n4563) );
  AOI22X1 U5455 ( .A(n2799), .B(inst_data_MEM_data[118]), .C(n4451), .D(
        inst_data_MEM_data[182]), .Y(n4562) );
  AND2X2 U5456 ( .A(n4563), .B(n4562), .Y(n4564) );
  NAND3X1 U5457 ( .A(n4566), .B(n4565), .C(n4564), .Y(u_MEM2WB_reg_N29) );
  AOI22X1 U5458 ( .A(n4609), .B(inst_data_MEM_data[23]), .C(n2800), .D(
        inst_data_MEM_data[215]), .Y(n4571) );
  AOI22X1 U5459 ( .A(n4437), .B(inst_data_MEM_data[55]), .C(n4451), .D(
        inst_data_MEM_data[183]), .Y(n4570) );
  AOI22X1 U5460 ( .A(n2798), .B(inst_data_MEM_data[151]), .C(n2797), .D(
        inst_data_MEM_data[247]), .Y(n4568) );
  AOI22X1 U5461 ( .A(n2799), .B(inst_data_MEM_data[119]), .C(n4602), .D(
        inst_data_MEM_data[87]), .Y(n4567) );
  AND2X2 U5462 ( .A(n4568), .B(n4567), .Y(n4569) );
  NAND3X1 U5463 ( .A(n4571), .B(n4570), .C(n4569), .Y(u_MEM2WB_reg_N30) );
  AOI22X1 U5464 ( .A(n2800), .B(inst_data_MEM_data[216]), .C(n4602), .D(
        inst_data_MEM_data[88]), .Y(n4576) );
  AOI22X1 U5465 ( .A(n4442), .B(inst_data_MEM_data[24]), .C(n4603), .D(
        inst_data_MEM_data[56]), .Y(n4575) );
  AOI22X1 U5466 ( .A(n2798), .B(inst_data_MEM_data[152]), .C(n4451), .D(
        inst_data_MEM_data[184]), .Y(n4573) );
  AOI22X1 U5467 ( .A(n2799), .B(inst_data_MEM_data[120]), .C(n2797), .D(
        inst_data_MEM_data[248]), .Y(n4572) );
  AND2X2 U5468 ( .A(n4573), .B(n4572), .Y(n4574) );
  NAND3X1 U5469 ( .A(n4576), .B(n4575), .C(n4574), .Y(u_MEM2WB_reg_N31) );
  AOI22X1 U5470 ( .A(n2799), .B(inst_data_MEM_data[121]), .C(n4451), .D(
        inst_data_MEM_data[185]), .Y(n4581) );
  AOI22X1 U5471 ( .A(n2798), .B(inst_data_MEM_data[153]), .C(n4602), .D(
        inst_data_MEM_data[89]), .Y(n4580) );
  AOI22X1 U5472 ( .A(n4609), .B(inst_data_MEM_data[25]), .C(n2800), .D(
        inst_data_MEM_data[217]), .Y(n4578) );
  AOI22X1 U5473 ( .A(n4437), .B(inst_data_MEM_data[57]), .C(n2797), .D(
        inst_data_MEM_data[249]), .Y(n4577) );
  AND2X2 U5474 ( .A(n4578), .B(n4577), .Y(n4579) );
  NAND3X1 U5475 ( .A(n4581), .B(n4580), .C(n4579), .Y(u_MEM2WB_reg_N32) );
  AOI22X1 U5476 ( .A(n4442), .B(inst_data_MEM_data[26]), .C(n2797), .D(
        inst_data_MEM_data[250]), .Y(n4586) );
  AOI22X1 U5477 ( .A(n4435), .B(inst_data_MEM_data[90]), .C(n4451), .D(
        inst_data_MEM_data[186]), .Y(n4585) );
  AOI22X1 U5478 ( .A(n2798), .B(inst_data_MEM_data[154]), .C(n2799), .D(
        inst_data_MEM_data[122]), .Y(n4583) );
  AOI22X1 U5479 ( .A(n2800), .B(inst_data_MEM_data[218]), .C(n4603), .D(
        inst_data_MEM_data[58]), .Y(n4582) );
  AND2X2 U5480 ( .A(n4583), .B(n4582), .Y(n4584) );
  NAND3X1 U5481 ( .A(n4586), .B(n4585), .C(n4584), .Y(u_MEM2WB_reg_N33) );
  AOI22X1 U5482 ( .A(n2798), .B(inst_data_MEM_data[155]), .C(n4435), .D(
        inst_data_MEM_data[91]), .Y(n4591) );
  AOI22X1 U5483 ( .A(n4442), .B(inst_data_MEM_data[27]), .C(n2797), .D(
        inst_data_MEM_data[251]), .Y(n4590) );
  AOI22X1 U5484 ( .A(n2800), .B(inst_data_MEM_data[219]), .C(n4437), .D(
        inst_data_MEM_data[59]), .Y(n4588) );
  AOI22X1 U5485 ( .A(n2799), .B(inst_data_MEM_data[123]), .C(n4451), .D(
        inst_data_MEM_data[187]), .Y(n4587) );
  AND2X2 U5486 ( .A(n4588), .B(n4587), .Y(n4589) );
  NAND3X1 U5487 ( .A(n4591), .B(n4590), .C(n4589), .Y(u_MEM2WB_reg_N34) );
  AOI22X1 U5488 ( .A(n2799), .B(inst_data_MEM_data[124]), .C(n2800), .D(
        inst_data_MEM_data[220]), .Y(n4596) );
  AOI22X1 U5489 ( .A(n2798), .B(inst_data_MEM_data[156]), .C(n4602), .D(
        inst_data_MEM_data[92]), .Y(n4595) );
  AOI22X1 U5490 ( .A(n4442), .B(inst_data_MEM_data[28]), .C(n4603), .D(
        inst_data_MEM_data[60]), .Y(n4593) );
  AOI22X1 U5491 ( .A(n4451), .B(inst_data_MEM_data[188]), .C(n2797), .D(
        inst_data_MEM_data[252]), .Y(n4592) );
  AND2X2 U5492 ( .A(n4593), .B(n4592), .Y(n4594) );
  NAND3X1 U5493 ( .A(n4596), .B(n4595), .C(n4594), .Y(u_MEM2WB_reg_N35) );
  AOI22X1 U5494 ( .A(n2799), .B(inst_data_MEM_data[125]), .C(n4435), .D(
        inst_data_MEM_data[93]), .Y(n4601) );
  AOI22X1 U5495 ( .A(n4437), .B(inst_data_MEM_data[61]), .C(n2797), .D(
        inst_data_MEM_data[253]), .Y(n4600) );
  AOI22X1 U5496 ( .A(n2800), .B(inst_data_MEM_data[221]), .C(n4451), .D(
        inst_data_MEM_data[189]), .Y(n4598) );
  AOI22X1 U5497 ( .A(n4442), .B(inst_data_MEM_data[29]), .C(n2798), .D(
        inst_data_MEM_data[157]), .Y(n4597) );
  AND2X2 U5498 ( .A(n4598), .B(n4597), .Y(n4599) );
  NAND3X1 U5499 ( .A(n4601), .B(n4600), .C(n4599), .Y(u_MEM2WB_reg_N36) );
  AOI22X1 U5500 ( .A(n4609), .B(inst_data_MEM_data[30]), .C(n2800), .D(
        inst_data_MEM_data[222]), .Y(n4608) );
  AOI22X1 U5501 ( .A(n2799), .B(inst_data_MEM_data[126]), .C(n4602), .D(
        inst_data_MEM_data[94]), .Y(n4607) );
  AOI22X1 U5502 ( .A(n4451), .B(inst_data_MEM_data[190]), .C(n2797), .D(
        inst_data_MEM_data[254]), .Y(n4605) );
  AOI22X1 U5503 ( .A(n2798), .B(inst_data_MEM_data[158]), .C(n4603), .D(
        inst_data_MEM_data[62]), .Y(n4604) );
  AND2X2 U5504 ( .A(n4605), .B(n4604), .Y(n4606) );
  NAND3X1 U5505 ( .A(n4608), .B(n4607), .C(n4606), .Y(u_MEM2WB_reg_N37) );
  AOI22X1 U5506 ( .A(n2800), .B(inst_data_MEM_data[223]), .C(n4437), .D(
        inst_data_MEM_data[63]), .Y(n4614) );
  AOI22X1 U5507 ( .A(n2799), .B(inst_data_MEM_data[127]), .C(n4451), .D(
        inst_data_MEM_data[191]), .Y(n4613) );
  AOI22X1 U5508 ( .A(n4609), .B(inst_data_MEM_data[31]), .C(n2797), .D(
        inst_data_MEM_data[255]), .Y(n4611) );
  AOI22X1 U5509 ( .A(n2798), .B(inst_data_MEM_data[159]), .C(n4435), .D(
        inst_data_MEM_data[95]), .Y(n4610) );
  AND2X2 U5510 ( .A(n4611), .B(n4610), .Y(n4612) );
  NAND3X1 U5511 ( .A(n4614), .B(n4613), .C(n4612), .Y(u_MEM2WB_reg_N38) );
  INVX1 U5512 ( .A(inst_address[30]), .Y(n4686) );
  INVX1 U5513 ( .A(inst_address[28]), .Y(n4691) );
  INVX1 U5514 ( .A(inst_address[26]), .Y(n4694) );
  NAND2X1 U5515 ( .A(inst_address[25]), .B(n4615), .Y(n5505) );
  NOR2X1 U5516 ( .A(n4694), .B(n5505), .Y(n5509) );
  NAND2X1 U5517 ( .A(inst_address[27]), .B(n5509), .Y(n5515) );
  NOR2X1 U5518 ( .A(n4691), .B(n5515), .Y(n5519) );
  INVX1 U5519 ( .A(inst_address[29]), .Y(n5522) );
  NOR2X1 U5520 ( .A(n5522), .B(n2796), .Y(n4687) );
  NAND3X1 U5521 ( .A(n4616), .B(n5519), .C(n4687), .Y(n5528) );
  AOI22X1 U5522 ( .A(n4617), .B(inst_address[31]), .C(n5526), .D(
        shifted_address_MEM[31]), .Y(n4618) );
  OAI21X1 U5523 ( .A(n4686), .B(n5528), .C(n4618), .Y(n2791) );
  INVX1 U5524 ( .A(instruction_ID[31]), .Y(n4620) );
  NAND2X1 U5525 ( .A(n4705), .B(instruction[31]), .Y(n4619) );
  OAI21X1 U5526 ( .A(n4620), .B(n5501), .C(n4619), .Y(n2790) );
  NAND2X1 U5527 ( .A(n4705), .B(instruction[30]), .Y(n4621) );
  OAI21X1 U5528 ( .A(n4622), .B(n5501), .C(n4621), .Y(n2789) );
  NAND2X1 U5529 ( .A(n4705), .B(instruction[29]), .Y(n4623) );
  OAI21X1 U5530 ( .A(n4624), .B(n4727), .C(n4623), .Y(n2788) );
  NAND2X1 U5531 ( .A(n4705), .B(instruction[28]), .Y(n4625) );
  OAI21X1 U5532 ( .A(n4626), .B(n4727), .C(n4625), .Y(n2787) );
  INVX1 U5533 ( .A(instruction_ID[27]), .Y(n4628) );
  NAND2X1 U5534 ( .A(n4705), .B(instruction[27]), .Y(n4627) );
  OAI21X1 U5535 ( .A(n4628), .B(n4727), .C(n4627), .Y(n2786) );
  INVX1 U5536 ( .A(instruction_ID[26]), .Y(n4630) );
  NAND2X1 U5537 ( .A(n4705), .B(instruction[26]), .Y(n4629) );
  OAI21X1 U5538 ( .A(n4630), .B(n5501), .C(n4629), .Y(n2785) );
  NAND2X1 U5539 ( .A(n4705), .B(instruction[25]), .Y(n4631) );
  OAI21X1 U5540 ( .A(n4727), .B(n4632), .C(n4631), .Y(n2784) );
  NAND2X1 U5541 ( .A(n4705), .B(instruction[24]), .Y(n4633) );
  OAI21X1 U5542 ( .A(n4727), .B(n4634), .C(n4633), .Y(n2783) );
  NAND2X1 U5543 ( .A(n4705), .B(instruction[23]), .Y(n4635) );
  OAI21X1 U5544 ( .A(n4727), .B(n4636), .C(n4635), .Y(n2782) );
  NAND2X1 U5545 ( .A(n4705), .B(instruction[22]), .Y(n4637) );
  OAI21X1 U5546 ( .A(n4727), .B(n4638), .C(n4637), .Y(n2781) );
  NAND2X1 U5547 ( .A(n4705), .B(instruction[21]), .Y(n4639) );
  OAI21X1 U5548 ( .A(n4727), .B(n4640), .C(n4639), .Y(n2780) );
  NAND2X1 U5549 ( .A(n4705), .B(instruction[20]), .Y(n4641) );
  OAI21X1 U5550 ( .A(n4727), .B(n4642), .C(n4641), .Y(n2779) );
  NAND2X1 U5551 ( .A(n4705), .B(instruction[19]), .Y(n4643) );
  OAI21X1 U5552 ( .A(n4727), .B(n4644), .C(n4643), .Y(n2778) );
  NAND2X1 U5553 ( .A(n4705), .B(instruction[18]), .Y(n4645) );
  OAI21X1 U5554 ( .A(n4727), .B(n4646), .C(n4645), .Y(n2777) );
  NAND2X1 U5555 ( .A(n4705), .B(instruction[17]), .Y(n4647) );
  OAI21X1 U5556 ( .A(n4727), .B(n4648), .C(n4647), .Y(n2776) );
  NAND2X1 U5557 ( .A(n4705), .B(instruction[16]), .Y(n4649) );
  OAI21X1 U5558 ( .A(n4727), .B(n4650), .C(n4649), .Y(n2775) );
  NAND2X1 U5559 ( .A(n4705), .B(instruction[15]), .Y(n4651) );
  OAI21X1 U5560 ( .A(n4652), .B(n5501), .C(n4651), .Y(n2774) );
  NAND2X1 U5561 ( .A(n4705), .B(instruction[14]), .Y(n4653) );
  OAI21X1 U5562 ( .A(n4654), .B(n4727), .C(n4653), .Y(n2773) );
  NAND2X1 U5563 ( .A(n4705), .B(instruction[13]), .Y(n4655) );
  OAI21X1 U5564 ( .A(n4656), .B(n5501), .C(n4655), .Y(n2772) );
  NAND2X1 U5565 ( .A(n4705), .B(instruction[12]), .Y(n4657) );
  OAI21X1 U5566 ( .A(n4658), .B(n4727), .C(n4657), .Y(n2771) );
  NAND2X1 U5567 ( .A(n4705), .B(instruction[11]), .Y(n4659) );
  OAI21X1 U5568 ( .A(n4660), .B(n5501), .C(n4659), .Y(n2770) );
  NAND2X1 U5569 ( .A(n4705), .B(instruction[10]), .Y(n4661) );
  OAI21X1 U5570 ( .A(n4662), .B(n5501), .C(n4661), .Y(n2769) );
  NAND2X1 U5571 ( .A(n4705), .B(instruction[9]), .Y(n4663) );
  OAI21X1 U5572 ( .A(n4664), .B(n4727), .C(n4663), .Y(n2768) );
  NAND2X1 U5573 ( .A(n4705), .B(instruction[8]), .Y(n4665) );
  OAI21X1 U5574 ( .A(n4666), .B(n4727), .C(n4665), .Y(n2767) );
  NAND2X1 U5575 ( .A(n4705), .B(instruction[7]), .Y(n4667) );
  OAI21X1 U5576 ( .A(n4668), .B(n5501), .C(n4667), .Y(n2766) );
  NAND2X1 U5577 ( .A(n4705), .B(instruction[6]), .Y(n4669) );
  OAI21X1 U5578 ( .A(n4670), .B(n5501), .C(n4669), .Y(n2765) );
  NAND2X1 U5579 ( .A(n4705), .B(instruction[5]), .Y(n4671) );
  OAI21X1 U5580 ( .A(n4672), .B(n4727), .C(n4671), .Y(n2764) );
  NAND2X1 U5581 ( .A(n4705), .B(instruction[4]), .Y(n4673) );
  OAI21X1 U5582 ( .A(n4674), .B(n5501), .C(n4673), .Y(n2763) );
  NAND2X1 U5583 ( .A(n4705), .B(instruction[3]), .Y(n4675) );
  OAI21X1 U5584 ( .A(n4676), .B(n5501), .C(n4675), .Y(n2762) );
  NAND2X1 U5585 ( .A(n4705), .B(instruction[2]), .Y(n4677) );
  OAI21X1 U5586 ( .A(n4678), .B(n4727), .C(n4677), .Y(n2761) );
  NAND2X1 U5587 ( .A(n4705), .B(instruction[1]), .Y(n4679) );
  OAI21X1 U5588 ( .A(n4680), .B(n5501), .C(n4679), .Y(n2760) );
  NAND2X1 U5589 ( .A(n4705), .B(instruction[0]), .Y(n4681) );
  OAI21X1 U5590 ( .A(n4682), .B(n5501), .C(n4681), .Y(n2759) );
  INVX1 U5591 ( .A(inst_address[31]), .Y(n4684) );
  OAI22X1 U5592 ( .A(n2796), .B(n4684), .C(n4727), .D(n4683), .Y(n2758) );
  OAI22X1 U5593 ( .A(n2796), .B(n4686), .C(n4727), .D(n4685), .Y(n2757) );
  OAI21X1 U5594 ( .A(n4727), .B(n4689), .C(n4688), .Y(n2756) );
  OAI22X1 U5595 ( .A(n2796), .B(n4691), .C(n4727), .D(n4690), .Y(n2755) );
  INVX1 U5596 ( .A(inst_address[27]), .Y(n5512) );
  OAI22X1 U5597 ( .A(n2796), .B(n5512), .C(n4727), .D(n4692), .Y(n2754) );
  OAI22X1 U5598 ( .A(n2796), .B(n4694), .C(n4727), .D(n4693), .Y(n2753) );
  INVX1 U5599 ( .A(inst_address[25]), .Y(n4696) );
  OAI22X1 U5600 ( .A(n2796), .B(n4696), .C(n4727), .D(n4695), .Y(n2752) );
  OAI22X1 U5601 ( .A(n2796), .B(n4698), .C(n5501), .D(n4697), .Y(n2751) );
  INVX1 U5602 ( .A(inst_address[23]), .Y(n4700) );
  OAI22X1 U5603 ( .A(n2796), .B(n4700), .C(n4727), .D(n4699), .Y(n2750) );
  OAI22X1 U5604 ( .A(n2796), .B(n4702), .C(n4727), .D(n4701), .Y(n2749) );
  INVX1 U5605 ( .A(inst_address[21]), .Y(n4704) );
  OAI22X1 U5606 ( .A(n2796), .B(n4704), .C(n4727), .D(n4703), .Y(n2748) );
  OAI22X1 U5607 ( .A(n2796), .B(n4707), .C(n4727), .D(n4706), .Y(n2747) );
  INVX1 U5608 ( .A(inst_address[19]), .Y(n4709) );
  OAI22X1 U5609 ( .A(n2796), .B(n4709), .C(n4727), .D(n4708), .Y(n2746) );
  OAI22X1 U5610 ( .A(n2796), .B(n4711), .C(n4727), .D(n4710), .Y(n2745) );
  OAI22X1 U5611 ( .A(n2796), .B(n4713), .C(n4727), .D(n4712), .Y(n2744) );
  INVX1 U5612 ( .A(inst_address[16]), .Y(n4715) );
  OAI22X1 U5613 ( .A(n2796), .B(n4715), .C(n4727), .D(n4714), .Y(n2743) );
  OAI22X1 U5614 ( .A(n2796), .B(n4717), .C(n4727), .D(n4716), .Y(n2742) );
  OAI22X1 U5615 ( .A(n2796), .B(n4719), .C(n4727), .D(n4718), .Y(n2741) );
  INVX1 U5616 ( .A(inst_address[13]), .Y(n4721) );
  OAI22X1 U5617 ( .A(n2796), .B(n4721), .C(n4727), .D(n4720), .Y(n2740) );
  OAI22X1 U5618 ( .A(n2796), .B(n4723), .C(n5501), .D(n4722), .Y(n2739) );
  INVX1 U5619 ( .A(inst_address[11]), .Y(n4725) );
  OAI22X1 U5620 ( .A(n2796), .B(n4725), .C(n5501), .D(n4724), .Y(n2738) );
  OAI22X1 U5621 ( .A(n2796), .B(n4728), .C(n4727), .D(n4726), .Y(n2737) );
  OAI22X1 U5622 ( .A(n2796), .B(n4730), .C(n5501), .D(n4729), .Y(n2736) );
  OAI22X1 U5623 ( .A(n2796), .B(n4732), .C(n5501), .D(n4731), .Y(n2735) );
  OAI22X1 U5624 ( .A(n2796), .B(n4734), .C(n5501), .D(n4733), .Y(n2734) );
  OAI22X1 U5625 ( .A(n2796), .B(n4736), .C(n5501), .D(n4735), .Y(n2733) );
  OAI22X1 U5626 ( .A(n2796), .B(n4738), .C(n5501), .D(n4737), .Y(n2732) );
  OAI22X1 U5627 ( .A(n2796), .B(n4740), .C(n5501), .D(n4739), .Y(n2731) );
  OAI22X1 U5628 ( .A(n2796), .B(n4742), .C(n5501), .D(n4741), .Y(n2730) );
  OAI22X1 U5629 ( .A(n2796), .B(n5502), .C(n5501), .D(n4743), .Y(n2729) );
  OAI22X1 U5630 ( .A(n2796), .B(n4745), .C(n5501), .D(n4744), .Y(n2728) );
  OAI22X1 U5631 ( .A(n2796), .B(n4747), .C(n5501), .D(n4746), .Y(n2727) );
  INVX1 U5632 ( .A(inst_data_MEM_data[255]), .Y(n4749) );
  INVX2 U5633 ( .A(n5014), .Y(n5062) );
  NAND2X1 U5634 ( .A(write_mem_data_MEM[31]), .B(n5062), .Y(n4748) );
  OAI21X1 U5635 ( .A(n5061), .B(n4749), .C(n4748), .Y(n2726) );
  NOR2X1 U5636 ( .A(write_mem_data_MEM[2]), .B(n5392), .Y(n4937) );
  AND2X2 U5637 ( .A(n4751), .B(n4927), .Y(n4753) );
  OAI21X1 U5638 ( .A(n5392), .B(inst_data_MEM_data[98]), .C(n5002), .Y(n4752)
         );
  OAI21X1 U5639 ( .A(n4937), .B(n5002), .C(n4752), .Y(n2725) );
  NAND2X1 U5640 ( .A(n2815), .B(write_mem_data_MEM[0]), .Y(n4891) );
  NOR2X1 U5641 ( .A(n4753), .B(n5392), .Y(n5000) );
  NAND2X1 U5642 ( .A(inst_data_MEM_data[96]), .B(n4754), .Y(n4755) );
  OAI21X1 U5643 ( .A(n4891), .B(n5002), .C(n4755), .Y(n2724) );
  NAND2X1 U5644 ( .A(n2815), .B(write_mem_data_MEM[1]), .Y(n4935) );
  NAND2X1 U5645 ( .A(inst_data_MEM_data[97]), .B(n4754), .Y(n4756) );
  OAI21X1 U5646 ( .A(n4935), .B(n5002), .C(n4756), .Y(n2723) );
  AND2X2 U5647 ( .A(n4758), .B(n4927), .Y(n4759) );
  NAND2X1 U5648 ( .A(n2815), .B(write_mem_data_MEM[31]), .Y(n5067) );
  NOR2X1 U5649 ( .A(n4759), .B(n5392), .Y(n4792) );
  NAND2X1 U5650 ( .A(inst_data_MEM_data[95]), .B(n4760), .Y(n4761) );
  OAI21X1 U5651 ( .A(n4794), .B(n5067), .C(n4761), .Y(n2722) );
  NOR2X1 U5652 ( .A(write_mem_data_MEM[0]), .B(n5392), .Y(n4933) );
  OAI21X1 U5653 ( .A(n5392), .B(inst_data_MEM_data[64]), .C(n4794), .Y(n4762)
         );
  OAI21X1 U5654 ( .A(n4933), .B(n4794), .C(n4762), .Y(n2721) );
  NOR2X1 U5655 ( .A(write_mem_data_MEM[1]), .B(n5392), .Y(n4893) );
  OAI21X1 U5656 ( .A(n5392), .B(inst_data_MEM_data[65]), .C(n4794), .Y(n4763)
         );
  OAI21X1 U5657 ( .A(n4893), .B(n4794), .C(n4763), .Y(n2720) );
  NAND2X1 U5658 ( .A(n2815), .B(write_mem_data_MEM[2]), .Y(n4841) );
  NAND2X1 U5659 ( .A(inst_data_MEM_data[66]), .B(n4760), .Y(n4764) );
  OAI21X1 U5660 ( .A(n4841), .B(n4794), .C(n4764), .Y(n2719) );
  NAND2X1 U5661 ( .A(n2815), .B(write_mem_data_MEM[3]), .Y(n4971) );
  NAND2X1 U5662 ( .A(inst_data_MEM_data[67]), .B(n4760), .Y(n4765) );
  OAI21X1 U5663 ( .A(n4971), .B(n4794), .C(n4765), .Y(n2718) );
  NAND2X1 U5664 ( .A(n2815), .B(write_mem_data_MEM[4]), .Y(n4973) );
  NAND2X1 U5665 ( .A(inst_data_MEM_data[68]), .B(n4760), .Y(n4766) );
  OAI21X1 U5666 ( .A(n4973), .B(n4794), .C(n4766), .Y(n2717) );
  NAND2X1 U5667 ( .A(n2815), .B(write_mem_data_MEM[5]), .Y(n4975) );
  NAND2X1 U5668 ( .A(inst_data_MEM_data[69]), .B(n4760), .Y(n4767) );
  OAI21X1 U5669 ( .A(n4975), .B(n4794), .C(n4767), .Y(n2716) );
  NAND2X1 U5670 ( .A(n2815), .B(write_mem_data_MEM[6]), .Y(n5069) );
  NAND2X1 U5671 ( .A(inst_data_MEM_data[70]), .B(n4760), .Y(n4768) );
  OAI21X1 U5672 ( .A(n5069), .B(n4794), .C(n4768), .Y(n2715) );
  NAND2X1 U5673 ( .A(n2815), .B(write_mem_data_MEM[7]), .Y(n5071) );
  NAND2X1 U5674 ( .A(inst_data_MEM_data[71]), .B(n4760), .Y(n4769) );
  OAI21X1 U5675 ( .A(n5071), .B(n4794), .C(n4769), .Y(n2714) );
  NAND2X1 U5676 ( .A(n2815), .B(write_mem_data_MEM[8]), .Y(n5073) );
  NAND2X1 U5677 ( .A(inst_data_MEM_data[72]), .B(n4760), .Y(n4770) );
  OAI21X1 U5678 ( .A(n5073), .B(n4794), .C(n4770), .Y(n2713) );
  NAND2X1 U5679 ( .A(n2815), .B(write_mem_data_MEM[9]), .Y(n5075) );
  NAND2X1 U5680 ( .A(inst_data_MEM_data[73]), .B(n4760), .Y(n4771) );
  OAI21X1 U5681 ( .A(n5075), .B(n4794), .C(n4771), .Y(n2712) );
  NAND2X1 U5682 ( .A(n3066), .B(write_mem_data_MEM[10]), .Y(n5077) );
  NAND2X1 U5683 ( .A(inst_data_MEM_data[74]), .B(n4760), .Y(n4772) );
  OAI21X1 U5684 ( .A(n5077), .B(n4794), .C(n4772), .Y(n2711) );
  NAND2X1 U5685 ( .A(n3066), .B(write_mem_data_MEM[11]), .Y(n5079) );
  NAND2X1 U5686 ( .A(inst_data_MEM_data[75]), .B(n4760), .Y(n4773) );
  OAI21X1 U5687 ( .A(n5079), .B(n4794), .C(n4773), .Y(n2710) );
  NAND2X1 U5688 ( .A(n3066), .B(write_mem_data_MEM[12]), .Y(n5081) );
  NAND2X1 U5689 ( .A(inst_data_MEM_data[76]), .B(n4760), .Y(n4774) );
  OAI21X1 U5690 ( .A(n5081), .B(n4794), .C(n4774), .Y(n2709) );
  NAND2X1 U5691 ( .A(n3066), .B(write_mem_data_MEM[13]), .Y(n5083) );
  NAND2X1 U5692 ( .A(inst_data_MEM_data[77]), .B(n4792), .Y(n4775) );
  OAI21X1 U5693 ( .A(n5083), .B(n4794), .C(n4775), .Y(n2708) );
  NAND2X1 U5694 ( .A(n3066), .B(write_mem_data_MEM[14]), .Y(n5085) );
  NAND2X1 U5695 ( .A(inst_data_MEM_data[78]), .B(n4792), .Y(n4776) );
  OAI21X1 U5696 ( .A(n5085), .B(n4794), .C(n4776), .Y(n2707) );
  NAND2X1 U5697 ( .A(n3066), .B(write_mem_data_MEM[15]), .Y(n5087) );
  NAND2X1 U5698 ( .A(inst_data_MEM_data[79]), .B(n4792), .Y(n4777) );
  OAI21X1 U5699 ( .A(n5087), .B(n4794), .C(n4777), .Y(n2706) );
  NAND2X1 U5700 ( .A(n3066), .B(write_mem_data_MEM[16]), .Y(n5089) );
  NAND2X1 U5701 ( .A(inst_data_MEM_data[80]), .B(n4760), .Y(n4778) );
  OAI21X1 U5702 ( .A(n5089), .B(n4794), .C(n4778), .Y(n2705) );
  NAND2X1 U5703 ( .A(n3066), .B(write_mem_data_MEM[17]), .Y(n5091) );
  NAND2X1 U5704 ( .A(inst_data_MEM_data[81]), .B(n4760), .Y(n4779) );
  OAI21X1 U5705 ( .A(n5091), .B(n4794), .C(n4779), .Y(n2704) );
  NAND2X1 U5706 ( .A(n3066), .B(write_mem_data_MEM[18]), .Y(n5093) );
  NAND2X1 U5707 ( .A(inst_data_MEM_data[82]), .B(n4792), .Y(n4780) );
  OAI21X1 U5708 ( .A(n5093), .B(n4794), .C(n4780), .Y(n2703) );
  NAND2X1 U5709 ( .A(n3066), .B(write_mem_data_MEM[19]), .Y(n5095) );
  NAND2X1 U5710 ( .A(inst_data_MEM_data[83]), .B(n4760), .Y(n4781) );
  OAI21X1 U5711 ( .A(n5095), .B(n4794), .C(n4781), .Y(n2702) );
  NAND2X1 U5712 ( .A(n3066), .B(write_mem_data_MEM[20]), .Y(n5097) );
  NAND2X1 U5713 ( .A(inst_data_MEM_data[84]), .B(n4760), .Y(n4782) );
  OAI21X1 U5714 ( .A(n5097), .B(n4794), .C(n4782), .Y(n2701) );
  NAND2X1 U5715 ( .A(n3066), .B(write_mem_data_MEM[21]), .Y(n5099) );
  NAND2X1 U5716 ( .A(inst_data_MEM_data[85]), .B(n4760), .Y(n4783) );
  OAI21X1 U5717 ( .A(n5099), .B(n4794), .C(n4783), .Y(n2700) );
  NAND2X1 U5718 ( .A(n3066), .B(write_mem_data_MEM[22]), .Y(n5101) );
  NAND2X1 U5719 ( .A(inst_data_MEM_data[86]), .B(n4760), .Y(n4784) );
  OAI21X1 U5720 ( .A(n5101), .B(n4794), .C(n4784), .Y(n2699) );
  NAND2X1 U5721 ( .A(n3066), .B(write_mem_data_MEM[23]), .Y(n5103) );
  NAND2X1 U5722 ( .A(inst_data_MEM_data[87]), .B(n4760), .Y(n4785) );
  OAI21X1 U5723 ( .A(n5103), .B(n4794), .C(n4785), .Y(n2698) );
  NAND2X1 U5724 ( .A(n3066), .B(write_mem_data_MEM[24]), .Y(n5105) );
  NAND2X1 U5725 ( .A(inst_data_MEM_data[88]), .B(n4760), .Y(n4786) );
  OAI21X1 U5726 ( .A(n5105), .B(n4794), .C(n4786), .Y(n2697) );
  NAND2X1 U5727 ( .A(n3066), .B(write_mem_data_MEM[25]), .Y(n5107) );
  NAND2X1 U5728 ( .A(inst_data_MEM_data[89]), .B(n4792), .Y(n4787) );
  OAI21X1 U5729 ( .A(n5107), .B(n4794), .C(n4787), .Y(n2696) );
  NAND2X1 U5730 ( .A(n3066), .B(write_mem_data_MEM[26]), .Y(n5109) );
  NAND2X1 U5731 ( .A(inst_data_MEM_data[90]), .B(n4792), .Y(n4788) );
  OAI21X1 U5732 ( .A(n5109), .B(n4794), .C(n4788), .Y(n2695) );
  NAND2X1 U5733 ( .A(n3066), .B(write_mem_data_MEM[27]), .Y(n5111) );
  NAND2X1 U5734 ( .A(inst_data_MEM_data[91]), .B(n4792), .Y(n4789) );
  OAI21X1 U5735 ( .A(n5111), .B(n4794), .C(n4789), .Y(n2694) );
  NAND2X1 U5736 ( .A(n3066), .B(write_mem_data_MEM[28]), .Y(n5114) );
  NAND2X1 U5737 ( .A(inst_data_MEM_data[92]), .B(n4792), .Y(n4790) );
  OAI21X1 U5738 ( .A(n5114), .B(n4794), .C(n4790), .Y(n2693) );
  NAND2X1 U5739 ( .A(n3066), .B(write_mem_data_MEM[29]), .Y(n5116) );
  NAND2X1 U5740 ( .A(inst_data_MEM_data[93]), .B(n4792), .Y(n4791) );
  OAI21X1 U5741 ( .A(n5116), .B(n4794), .C(n4791), .Y(n2692) );
  NAND2X1 U5742 ( .A(n3066), .B(write_mem_data_MEM[30]), .Y(n5118) );
  NAND2X1 U5743 ( .A(inst_data_MEM_data[94]), .B(n4792), .Y(n4793) );
  OAI21X1 U5744 ( .A(n5118), .B(n4794), .C(n4793), .Y(n2691) );
  NAND2X1 U5745 ( .A(n4795), .B(n4927), .Y(n4832) );
  INVX2 U5746 ( .A(n4796), .Y(n4829) );
  NOR2X1 U5747 ( .A(n4796), .B(n5392), .Y(n4830) );
  NAND2X1 U5748 ( .A(inst_data_MEM_data[63]), .B(n4797), .Y(n4798) );
  OAI21X1 U5749 ( .A(n4829), .B(n5067), .C(n4798), .Y(n2690) );
  NAND2X1 U5750 ( .A(inst_data_MEM_data[32]), .B(n4797), .Y(n4799) );
  OAI21X1 U5751 ( .A(n4829), .B(n4891), .C(n4799), .Y(n2689) );
  OAI21X1 U5752 ( .A(n5392), .B(inst_data_MEM_data[33]), .C(n4829), .Y(n4800)
         );
  OAI21X1 U5753 ( .A(n4893), .B(n4829), .C(n4800), .Y(n2688) );
  NAND2X1 U5754 ( .A(inst_data_MEM_data[34]), .B(n4797), .Y(n4801) );
  OAI21X1 U5755 ( .A(n4829), .B(n4841), .C(n4801), .Y(n2687) );
  NAND2X1 U5756 ( .A(inst_data_MEM_data[35]), .B(n4797), .Y(n4802) );
  OAI21X1 U5757 ( .A(n4829), .B(n4971), .C(n4802), .Y(n2686) );
  NAND2X1 U5758 ( .A(inst_data_MEM_data[36]), .B(n4797), .Y(n4803) );
  OAI21X1 U5759 ( .A(n4829), .B(n4973), .C(n4803), .Y(n2685) );
  NAND2X1 U5760 ( .A(inst_data_MEM_data[37]), .B(n4797), .Y(n4804) );
  OAI21X1 U5761 ( .A(n4829), .B(n4975), .C(n4804), .Y(n2684) );
  NAND2X1 U5762 ( .A(inst_data_MEM_data[38]), .B(n4797), .Y(n4805) );
  OAI21X1 U5763 ( .A(n4829), .B(n5069), .C(n4805), .Y(n2683) );
  NAND2X1 U5764 ( .A(inst_data_MEM_data[39]), .B(n4797), .Y(n4806) );
  OAI21X1 U5765 ( .A(n4832), .B(n5071), .C(n4806), .Y(n2682) );
  NAND2X1 U5766 ( .A(inst_data_MEM_data[40]), .B(n4797), .Y(n4807) );
  OAI21X1 U5767 ( .A(n4832), .B(n5073), .C(n4807), .Y(n2681) );
  NAND2X1 U5768 ( .A(inst_data_MEM_data[41]), .B(n4797), .Y(n4808) );
  OAI21X1 U5769 ( .A(n4832), .B(n5075), .C(n4808), .Y(n2680) );
  NAND2X1 U5770 ( .A(inst_data_MEM_data[42]), .B(n4797), .Y(n4809) );
  OAI21X1 U5771 ( .A(n4832), .B(n5077), .C(n4809), .Y(n2679) );
  NAND2X1 U5772 ( .A(inst_data_MEM_data[43]), .B(n4797), .Y(n4810) );
  OAI21X1 U5773 ( .A(n4832), .B(n5079), .C(n4810), .Y(n2678) );
  NAND2X1 U5774 ( .A(inst_data_MEM_data[44]), .B(n4830), .Y(n4811) );
  OAI21X1 U5775 ( .A(n4832), .B(n5081), .C(n4811), .Y(n2677) );
  NAND2X1 U5776 ( .A(inst_data_MEM_data[45]), .B(n4830), .Y(n4812) );
  OAI21X1 U5777 ( .A(n4832), .B(n5083), .C(n4812), .Y(n2676) );
  NAND2X1 U5778 ( .A(inst_data_MEM_data[46]), .B(n4830), .Y(n4813) );
  OAI21X1 U5779 ( .A(n4832), .B(n5085), .C(n4813), .Y(n2675) );
  NAND2X1 U5780 ( .A(inst_data_MEM_data[47]), .B(n4830), .Y(n4814) );
  OAI21X1 U5781 ( .A(n4832), .B(n5087), .C(n4814), .Y(n2674) );
  NAND2X1 U5782 ( .A(inst_data_MEM_data[48]), .B(n4830), .Y(n4815) );
  OAI21X1 U5783 ( .A(n4832), .B(n5089), .C(n4815), .Y(n2673) );
  NAND2X1 U5784 ( .A(inst_data_MEM_data[49]), .B(n4830), .Y(n4816) );
  OAI21X1 U5785 ( .A(n4829), .B(n5091), .C(n4816), .Y(n2672) );
  NAND2X1 U5786 ( .A(inst_data_MEM_data[50]), .B(n4830), .Y(n4817) );
  OAI21X1 U5787 ( .A(n4832), .B(n5093), .C(n4817), .Y(n2671) );
  NAND2X1 U5788 ( .A(inst_data_MEM_data[51]), .B(n4830), .Y(n4818) );
  OAI21X1 U5789 ( .A(n4829), .B(n5095), .C(n4818), .Y(n2670) );
  NAND2X1 U5790 ( .A(inst_data_MEM_data[52]), .B(n4797), .Y(n4819) );
  OAI21X1 U5791 ( .A(n4829), .B(n5097), .C(n4819), .Y(n2669) );
  NAND2X1 U5792 ( .A(inst_data_MEM_data[53]), .B(n4797), .Y(n4820) );
  OAI21X1 U5793 ( .A(n4829), .B(n5099), .C(n4820), .Y(n2668) );
  NAND2X1 U5794 ( .A(inst_data_MEM_data[54]), .B(n4830), .Y(n4821) );
  OAI21X1 U5795 ( .A(n4829), .B(n5101), .C(n4821), .Y(n2667) );
  NAND2X1 U5796 ( .A(inst_data_MEM_data[55]), .B(n4830), .Y(n4822) );
  OAI21X1 U5797 ( .A(n4829), .B(n5103), .C(n4822), .Y(n2666) );
  NAND2X1 U5798 ( .A(inst_data_MEM_data[56]), .B(n4830), .Y(n4823) );
  OAI21X1 U5799 ( .A(n4829), .B(n5105), .C(n4823), .Y(n2665) );
  NAND2X1 U5800 ( .A(inst_data_MEM_data[57]), .B(n4797), .Y(n4824) );
  OAI21X1 U5801 ( .A(n4829), .B(n5107), .C(n4824), .Y(n2664) );
  NAND2X1 U5802 ( .A(inst_data_MEM_data[58]), .B(n4830), .Y(n4825) );
  OAI21X1 U5803 ( .A(n4829), .B(n5109), .C(n4825), .Y(n2663) );
  NAND2X1 U5804 ( .A(inst_data_MEM_data[59]), .B(n4830), .Y(n4826) );
  OAI21X1 U5805 ( .A(n4829), .B(n5111), .C(n4826), .Y(n2662) );
  NAND2X1 U5806 ( .A(inst_data_MEM_data[60]), .B(n4830), .Y(n4827) );
  OAI21X1 U5807 ( .A(n4829), .B(n5114), .C(n4827), .Y(n2661) );
  NAND2X1 U5808 ( .A(inst_data_MEM_data[61]), .B(n4830), .Y(n4828) );
  OAI21X1 U5809 ( .A(n4829), .B(n5116), .C(n4828), .Y(n2660) );
  NAND2X1 U5810 ( .A(inst_data_MEM_data[62]), .B(n4830), .Y(n4831) );
  OAI21X1 U5811 ( .A(n4832), .B(n5118), .C(n4831), .Y(n2659) );
  NAND2X1 U5812 ( .A(n4834), .B(n4927), .Y(n4872) );
  INVX2 U5813 ( .A(n4835), .Y(n4869) );
  NOR2X1 U5814 ( .A(n4835), .B(n5392), .Y(n4870) );
  NAND2X1 U5815 ( .A(inst_data_MEM_data[31]), .B(n4836), .Y(n4837) );
  OAI21X1 U5816 ( .A(n4869), .B(n5067), .C(n4837), .Y(n2658) );
  OAI21X1 U5817 ( .A(n5392), .B(inst_data_MEM_data[0]), .C(n4869), .Y(n4838)
         );
  OAI21X1 U5818 ( .A(n4933), .B(n4869), .C(n4838), .Y(n2657) );
  NAND2X1 U5819 ( .A(inst_data_MEM_data[1]), .B(n4836), .Y(n4839) );
  OAI21X1 U5820 ( .A(n4869), .B(n4935), .C(n4839), .Y(n2656) );
  NAND2X1 U5821 ( .A(inst_data_MEM_data[2]), .B(n4836), .Y(n4840) );
  OAI21X1 U5822 ( .A(n4869), .B(n4841), .C(n4840), .Y(n2655) );
  NAND2X1 U5823 ( .A(inst_data_MEM_data[3]), .B(n4836), .Y(n4842) );
  OAI21X1 U5824 ( .A(n4869), .B(n4971), .C(n4842), .Y(n2654) );
  NAND2X1 U5825 ( .A(inst_data_MEM_data[4]), .B(n4836), .Y(n4843) );
  OAI21X1 U5826 ( .A(n4869), .B(n4973), .C(n4843), .Y(n2653) );
  NAND2X1 U5827 ( .A(inst_data_MEM_data[5]), .B(n4836), .Y(n4844) );
  OAI21X1 U5828 ( .A(n4869), .B(n4975), .C(n4844), .Y(n2652) );
  NAND2X1 U5829 ( .A(inst_data_MEM_data[6]), .B(n4836), .Y(n4845) );
  OAI21X1 U5830 ( .A(n4869), .B(n5069), .C(n4845), .Y(n2651) );
  NAND2X1 U5831 ( .A(inst_data_MEM_data[7]), .B(n4836), .Y(n4846) );
  OAI21X1 U5832 ( .A(n4872), .B(n5071), .C(n4846), .Y(n2650) );
  NAND2X1 U5833 ( .A(inst_data_MEM_data[8]), .B(n4836), .Y(n4847) );
  OAI21X1 U5834 ( .A(n4872), .B(n5073), .C(n4847), .Y(n2649) );
  NAND2X1 U5835 ( .A(inst_data_MEM_data[9]), .B(n4836), .Y(n4848) );
  OAI21X1 U5836 ( .A(n4872), .B(n5075), .C(n4848), .Y(n2648) );
  NAND2X1 U5837 ( .A(inst_data_MEM_data[10]), .B(n4836), .Y(n4849) );
  OAI21X1 U5838 ( .A(n4872), .B(n5077), .C(n4849), .Y(n2647) );
  NAND2X1 U5839 ( .A(inst_data_MEM_data[11]), .B(n4836), .Y(n4850) );
  OAI21X1 U5840 ( .A(n4872), .B(n5079), .C(n4850), .Y(n2646) );
  NAND2X1 U5841 ( .A(inst_data_MEM_data[12]), .B(n4870), .Y(n4851) );
  OAI21X1 U5842 ( .A(n4872), .B(n5081), .C(n4851), .Y(n2645) );
  NAND2X1 U5843 ( .A(inst_data_MEM_data[13]), .B(n4870), .Y(n4852) );
  OAI21X1 U5844 ( .A(n4872), .B(n5083), .C(n4852), .Y(n2644) );
  NAND2X1 U5845 ( .A(inst_data_MEM_data[14]), .B(n4870), .Y(n4853) );
  OAI21X1 U5846 ( .A(n4872), .B(n5085), .C(n4853), .Y(n2643) );
  NAND2X1 U5847 ( .A(inst_data_MEM_data[15]), .B(n4870), .Y(n4854) );
  OAI21X1 U5848 ( .A(n4872), .B(n5087), .C(n4854), .Y(n2642) );
  NAND2X1 U5849 ( .A(inst_data_MEM_data[16]), .B(n4870), .Y(n4855) );
  OAI21X1 U5850 ( .A(n4872), .B(n5089), .C(n4855), .Y(n2641) );
  NAND2X1 U5851 ( .A(inst_data_MEM_data[17]), .B(n4870), .Y(n4856) );
  OAI21X1 U5852 ( .A(n4869), .B(n5091), .C(n4856), .Y(n2640) );
  NAND2X1 U5853 ( .A(inst_data_MEM_data[18]), .B(n4870), .Y(n4857) );
  OAI21X1 U5854 ( .A(n4872), .B(n5093), .C(n4857), .Y(n2639) );
  NAND2X1 U5855 ( .A(inst_data_MEM_data[19]), .B(n4870), .Y(n4858) );
  OAI21X1 U5856 ( .A(n4869), .B(n5095), .C(n4858), .Y(n2638) );
  NAND2X1 U5857 ( .A(inst_data_MEM_data[20]), .B(n4870), .Y(n4859) );
  OAI21X1 U5858 ( .A(n4869), .B(n5097), .C(n4859), .Y(n2637) );
  NAND2X1 U5859 ( .A(inst_data_MEM_data[21]), .B(n4870), .Y(n4860) );
  OAI21X1 U5860 ( .A(n4869), .B(n5099), .C(n4860), .Y(n2636) );
  NAND2X1 U5861 ( .A(inst_data_MEM_data[22]), .B(n4836), .Y(n4861) );
  OAI21X1 U5862 ( .A(n4869), .B(n5101), .C(n4861), .Y(n2635) );
  NAND2X1 U5863 ( .A(inst_data_MEM_data[23]), .B(n4836), .Y(n4862) );
  OAI21X1 U5864 ( .A(n4869), .B(n5103), .C(n4862), .Y(n2634) );
  NAND2X1 U5865 ( .A(inst_data_MEM_data[24]), .B(n4836), .Y(n4863) );
  OAI21X1 U5866 ( .A(n4869), .B(n5105), .C(n4863), .Y(n2633) );
  NAND2X1 U5867 ( .A(inst_data_MEM_data[25]), .B(n4870), .Y(n4864) );
  OAI21X1 U5868 ( .A(n4869), .B(n5107), .C(n4864), .Y(n2632) );
  NAND2X1 U5869 ( .A(inst_data_MEM_data[26]), .B(n4870), .Y(n4865) );
  OAI21X1 U5870 ( .A(n4869), .B(n5109), .C(n4865), .Y(n2631) );
  NAND2X1 U5871 ( .A(inst_data_MEM_data[27]), .B(n4870), .Y(n4866) );
  OAI21X1 U5872 ( .A(n4869), .B(n5111), .C(n4866), .Y(n2630) );
  NAND2X1 U5873 ( .A(inst_data_MEM_data[28]), .B(n4870), .Y(n4867) );
  OAI21X1 U5874 ( .A(n4869), .B(n5114), .C(n4867), .Y(n2629) );
  NAND2X1 U5875 ( .A(inst_data_MEM_data[29]), .B(n4870), .Y(n4868) );
  OAI21X1 U5876 ( .A(n4869), .B(n5116), .C(n4868), .Y(n2628) );
  NAND2X1 U5877 ( .A(inst_data_MEM_data[30]), .B(n4870), .Y(n4871) );
  OAI21X1 U5878 ( .A(n4872), .B(n5118), .C(n4871), .Y(n2627) );
  INVX1 U5879 ( .A(inst_data_MEM_data[254]), .Y(n4874) );
  NAND2X1 U5880 ( .A(n5062), .B(write_mem_data_MEM[30]), .Y(n4873) );
  OAI21X1 U5881 ( .A(n5065), .B(n4874), .C(n4873), .Y(n2626) );
  AND2X2 U5882 ( .A(n4876), .B(n4927), .Y(n4877) );
  NOR2X1 U5883 ( .A(n4877), .B(n5392), .Y(n5112) );
  NAND2X1 U5884 ( .A(inst_data_MEM_data[197]), .B(n4878), .Y(n4879) );
  OAI21X1 U5885 ( .A(n5119), .B(n4975), .C(n4879), .Y(n2625) );
  OAI21X1 U5886 ( .A(n5392), .B(inst_data_MEM_data[192]), .C(n5119), .Y(n4880)
         );
  OAI21X1 U5887 ( .A(n4933), .B(n5119), .C(n4880), .Y(n2624) );
  OAI21X1 U5888 ( .A(n5392), .B(inst_data_MEM_data[193]), .C(n5119), .Y(n4881)
         );
  OAI21X1 U5889 ( .A(n4893), .B(n5119), .C(n4881), .Y(n2623) );
  OAI21X1 U5890 ( .A(n5392), .B(inst_data_MEM_data[194]), .C(n5119), .Y(n4882)
         );
  OAI21X1 U5891 ( .A(n4937), .B(n5119), .C(n4882), .Y(n2622) );
  NAND2X1 U5892 ( .A(inst_data_MEM_data[195]), .B(n4878), .Y(n4883) );
  OAI21X1 U5893 ( .A(n5119), .B(n4971), .C(n4883), .Y(n2621) );
  NAND2X1 U5894 ( .A(inst_data_MEM_data[196]), .B(n4878), .Y(n4884) );
  OAI21X1 U5895 ( .A(n5119), .B(n4973), .C(n4884), .Y(n2620) );
  NAND2X1 U5896 ( .A(n4886), .B(n4927), .Y(n4925) );
  NOR2X1 U5897 ( .A(n4889), .B(n5392), .Y(n4923) );
  NAND2X1 U5898 ( .A(inst_data_MEM_data[191]), .B(n4887), .Y(n4888) );
  OAI21X1 U5899 ( .A(n4925), .B(n5067), .C(n4888), .Y(n2619) );
  INVX2 U5900 ( .A(n4889), .Y(n4922) );
  NAND2X1 U5901 ( .A(inst_data_MEM_data[160]), .B(n4887), .Y(n4890) );
  OAI21X1 U5902 ( .A(n4922), .B(n4891), .C(n4890), .Y(n2618) );
  OAI21X1 U5903 ( .A(n5392), .B(inst_data_MEM_data[161]), .C(n4922), .Y(n4892)
         );
  OAI21X1 U5904 ( .A(n4893), .B(n4922), .C(n4892), .Y(n2617) );
  OAI21X1 U5905 ( .A(n5392), .B(inst_data_MEM_data[162]), .C(n4922), .Y(n4894)
         );
  OAI21X1 U5906 ( .A(n4937), .B(n4922), .C(n4894), .Y(n2616) );
  NAND2X1 U5907 ( .A(inst_data_MEM_data[163]), .B(n4887), .Y(n4895) );
  OAI21X1 U5908 ( .A(n4922), .B(n4971), .C(n4895), .Y(n2615) );
  NAND2X1 U5909 ( .A(inst_data_MEM_data[164]), .B(n4887), .Y(n4896) );
  OAI21X1 U5910 ( .A(n4922), .B(n4973), .C(n4896), .Y(n2614) );
  NAND2X1 U5911 ( .A(inst_data_MEM_data[165]), .B(n4887), .Y(n4897) );
  OAI21X1 U5912 ( .A(n4922), .B(n4975), .C(n4897), .Y(n2613) );
  NAND2X1 U5913 ( .A(inst_data_MEM_data[166]), .B(n4887), .Y(n4898) );
  OAI21X1 U5914 ( .A(n4922), .B(n5069), .C(n4898), .Y(n2612) );
  NAND2X1 U5915 ( .A(inst_data_MEM_data[167]), .B(n4887), .Y(n4899) );
  OAI21X1 U5916 ( .A(n4922), .B(n5071), .C(n4899), .Y(n2611) );
  NAND2X1 U5917 ( .A(inst_data_MEM_data[168]), .B(n4887), .Y(n4900) );
  OAI21X1 U5918 ( .A(n4925), .B(n5073), .C(n4900), .Y(n2610) );
  NAND2X1 U5919 ( .A(inst_data_MEM_data[169]), .B(n4887), .Y(n4901) );
  OAI21X1 U5920 ( .A(n4925), .B(n5075), .C(n4901), .Y(n2609) );
  NAND2X1 U5921 ( .A(inst_data_MEM_data[170]), .B(n4887), .Y(n4902) );
  OAI21X1 U5922 ( .A(n4925), .B(n5077), .C(n4902), .Y(n2608) );
  NAND2X1 U5923 ( .A(inst_data_MEM_data[171]), .B(n4887), .Y(n4903) );
  OAI21X1 U5924 ( .A(n4925), .B(n5079), .C(n4903), .Y(n2607) );
  NAND2X1 U5925 ( .A(inst_data_MEM_data[172]), .B(n4887), .Y(n4904) );
  OAI21X1 U5926 ( .A(n4925), .B(n5081), .C(n4904), .Y(n2606) );
  NAND2X1 U5927 ( .A(inst_data_MEM_data[173]), .B(n4923), .Y(n4905) );
  OAI21X1 U5928 ( .A(n4925), .B(n5083), .C(n4905), .Y(n2605) );
  NAND2X1 U5929 ( .A(inst_data_MEM_data[174]), .B(n4923), .Y(n4906) );
  OAI21X1 U5930 ( .A(n4925), .B(n5085), .C(n4906), .Y(n2604) );
  NAND2X1 U5931 ( .A(inst_data_MEM_data[175]), .B(n4923), .Y(n4907) );
  OAI21X1 U5932 ( .A(n4925), .B(n5087), .C(n4907), .Y(n2603) );
  NAND2X1 U5933 ( .A(inst_data_MEM_data[176]), .B(n4923), .Y(n4908) );
  OAI21X1 U5934 ( .A(n4925), .B(n5089), .C(n4908), .Y(n2602) );
  NAND2X1 U5935 ( .A(inst_data_MEM_data[177]), .B(n4887), .Y(n4909) );
  OAI21X1 U5936 ( .A(n4925), .B(n5091), .C(n4909), .Y(n2601) );
  NAND2X1 U5937 ( .A(inst_data_MEM_data[178]), .B(n4887), .Y(n4910) );
  OAI21X1 U5938 ( .A(n4922), .B(n5093), .C(n4910), .Y(n2600) );
  NAND2X1 U5939 ( .A(inst_data_MEM_data[179]), .B(n4887), .Y(n4911) );
  OAI21X1 U5940 ( .A(n4922), .B(n5095), .C(n4911), .Y(n2599) );
  NAND2X1 U5941 ( .A(inst_data_MEM_data[180]), .B(n4887), .Y(n4912) );
  OAI21X1 U5942 ( .A(n4922), .B(n5097), .C(n4912), .Y(n2598) );
  NAND2X1 U5943 ( .A(inst_data_MEM_data[181]), .B(n4887), .Y(n4913) );
  OAI21X1 U5944 ( .A(n4922), .B(n5099), .C(n4913), .Y(n2597) );
  NAND2X1 U5945 ( .A(inst_data_MEM_data[182]), .B(n4887), .Y(n4914) );
  OAI21X1 U5946 ( .A(n4922), .B(n5101), .C(n4914), .Y(n2596) );
  NAND2X1 U5947 ( .A(inst_data_MEM_data[183]), .B(n4887), .Y(n4915) );
  OAI21X1 U5948 ( .A(n4922), .B(n5103), .C(n4915), .Y(n2595) );
  NAND2X1 U5949 ( .A(inst_data_MEM_data[184]), .B(n4887), .Y(n4916) );
  OAI21X1 U5950 ( .A(n4922), .B(n5105), .C(n4916), .Y(n2594) );
  NAND2X1 U5951 ( .A(inst_data_MEM_data[185]), .B(n4923), .Y(n4917) );
  OAI21X1 U5952 ( .A(n4922), .B(n5107), .C(n4917), .Y(n2593) );
  NAND2X1 U5953 ( .A(inst_data_MEM_data[186]), .B(n4923), .Y(n4918) );
  OAI21X1 U5954 ( .A(n4922), .B(n5109), .C(n4918), .Y(n2592) );
  NAND2X1 U5955 ( .A(inst_data_MEM_data[187]), .B(n4923), .Y(n4919) );
  OAI21X1 U5956 ( .A(n4922), .B(n5111), .C(n4919), .Y(n2591) );
  NAND2X1 U5957 ( .A(inst_data_MEM_data[188]), .B(n4923), .Y(n4920) );
  OAI21X1 U5958 ( .A(n4922), .B(n5114), .C(n4920), .Y(n2590) );
  NAND2X1 U5959 ( .A(inst_data_MEM_data[189]), .B(n4923), .Y(n4921) );
  OAI21X1 U5960 ( .A(n4922), .B(n5116), .C(n4921), .Y(n2589) );
  NAND2X1 U5961 ( .A(inst_data_MEM_data[190]), .B(n4923), .Y(n4924) );
  OAI21X1 U5962 ( .A(n4925), .B(n5118), .C(n4924), .Y(n2588) );
  NAND2X1 U5963 ( .A(n4928), .B(n4927), .Y(n4968) );
  NOR2X1 U5964 ( .A(n4931), .B(n5392), .Y(n4966) );
  NAND2X1 U5965 ( .A(inst_data_MEM_data[159]), .B(n4929), .Y(n4930) );
  OAI21X1 U5966 ( .A(n4968), .B(n5067), .C(n4930), .Y(n2587) );
  INVX2 U5967 ( .A(n4931), .Y(n4965) );
  OAI21X1 U5968 ( .A(n5392), .B(inst_data_MEM_data[128]), .C(n4965), .Y(n4932)
         );
  OAI21X1 U5969 ( .A(n4933), .B(n4965), .C(n4932), .Y(n2586) );
  NAND2X1 U5970 ( .A(inst_data_MEM_data[129]), .B(n4929), .Y(n4934) );
  OAI21X1 U5971 ( .A(n4965), .B(n4935), .C(n4934), .Y(n2585) );
  OAI21X1 U5972 ( .A(n5392), .B(inst_data_MEM_data[130]), .C(n4965), .Y(n4936)
         );
  OAI21X1 U5973 ( .A(n4937), .B(n4965), .C(n4936), .Y(n2584) );
  NAND2X1 U5974 ( .A(inst_data_MEM_data[131]), .B(n4929), .Y(n4938) );
  OAI21X1 U5975 ( .A(n4965), .B(n4971), .C(n4938), .Y(n2583) );
  NAND2X1 U5976 ( .A(inst_data_MEM_data[132]), .B(n4929), .Y(n4939) );
  OAI21X1 U5977 ( .A(n4965), .B(n4973), .C(n4939), .Y(n2582) );
  NAND2X1 U5978 ( .A(inst_data_MEM_data[133]), .B(n4929), .Y(n4940) );
  OAI21X1 U5979 ( .A(n4965), .B(n4975), .C(n4940), .Y(n2581) );
  NAND2X1 U5980 ( .A(inst_data_MEM_data[134]), .B(n4929), .Y(n4941) );
  OAI21X1 U5981 ( .A(n4965), .B(n5069), .C(n4941), .Y(n2580) );
  NAND2X1 U5982 ( .A(inst_data_MEM_data[135]), .B(n4929), .Y(n4942) );
  OAI21X1 U5983 ( .A(n4965), .B(n5071), .C(n4942), .Y(n2579) );
  NAND2X1 U5984 ( .A(inst_data_MEM_data[136]), .B(n4929), .Y(n4943) );
  OAI21X1 U5985 ( .A(n4968), .B(n5073), .C(n4943), .Y(n2578) );
  NAND2X1 U5986 ( .A(inst_data_MEM_data[137]), .B(n4929), .Y(n4944) );
  OAI21X1 U5987 ( .A(n4968), .B(n5075), .C(n4944), .Y(n2577) );
  NAND2X1 U5988 ( .A(inst_data_MEM_data[138]), .B(n4929), .Y(n4945) );
  OAI21X1 U5989 ( .A(n4968), .B(n5077), .C(n4945), .Y(n2576) );
  NAND2X1 U5990 ( .A(inst_data_MEM_data[139]), .B(n4929), .Y(n4946) );
  OAI21X1 U5991 ( .A(n4968), .B(n5079), .C(n4946), .Y(n2575) );
  NAND2X1 U5992 ( .A(inst_data_MEM_data[140]), .B(n4929), .Y(n4947) );
  OAI21X1 U5993 ( .A(n4968), .B(n5081), .C(n4947), .Y(n2574) );
  NAND2X1 U5994 ( .A(inst_data_MEM_data[141]), .B(n4966), .Y(n4948) );
  OAI21X1 U5995 ( .A(n4968), .B(n5083), .C(n4948), .Y(n2573) );
  NAND2X1 U5996 ( .A(inst_data_MEM_data[142]), .B(n4966), .Y(n4949) );
  OAI21X1 U5997 ( .A(n4968), .B(n5085), .C(n4949), .Y(n2572) );
  NAND2X1 U5998 ( .A(inst_data_MEM_data[143]), .B(n4966), .Y(n4950) );
  OAI21X1 U5999 ( .A(n4968), .B(n5087), .C(n4950), .Y(n2571) );
  NAND2X1 U6000 ( .A(inst_data_MEM_data[144]), .B(n4966), .Y(n4951) );
  OAI21X1 U6001 ( .A(n4968), .B(n5089), .C(n4951), .Y(n2570) );
  NAND2X1 U6002 ( .A(inst_data_MEM_data[145]), .B(n4929), .Y(n4952) );
  OAI21X1 U6003 ( .A(n4968), .B(n5091), .C(n4952), .Y(n2569) );
  NAND2X1 U6004 ( .A(inst_data_MEM_data[146]), .B(n4929), .Y(n4953) );
  OAI21X1 U6005 ( .A(n4965), .B(n5093), .C(n4953), .Y(n2568) );
  NAND2X1 U6006 ( .A(inst_data_MEM_data[147]), .B(n4929), .Y(n4954) );
  OAI21X1 U6007 ( .A(n4965), .B(n5095), .C(n4954), .Y(n2567) );
  NAND2X1 U6008 ( .A(inst_data_MEM_data[148]), .B(n4929), .Y(n4955) );
  OAI21X1 U6009 ( .A(n4965), .B(n5097), .C(n4955), .Y(n2566) );
  NAND2X1 U6010 ( .A(inst_data_MEM_data[149]), .B(n4929), .Y(n4956) );
  OAI21X1 U6011 ( .A(n4965), .B(n5099), .C(n4956), .Y(n2565) );
  NAND2X1 U6012 ( .A(inst_data_MEM_data[150]), .B(n4929), .Y(n4957) );
  OAI21X1 U6013 ( .A(n4965), .B(n5101), .C(n4957), .Y(n2564) );
  NAND2X1 U6014 ( .A(inst_data_MEM_data[151]), .B(n4929), .Y(n4958) );
  OAI21X1 U6015 ( .A(n4965), .B(n5103), .C(n4958), .Y(n2563) );
  NAND2X1 U6016 ( .A(inst_data_MEM_data[152]), .B(n4929), .Y(n4959) );
  OAI21X1 U6017 ( .A(n4965), .B(n5105), .C(n4959), .Y(n2562) );
  NAND2X1 U6018 ( .A(inst_data_MEM_data[153]), .B(n4966), .Y(n4960) );
  OAI21X1 U6019 ( .A(n4965), .B(n5107), .C(n4960), .Y(n2561) );
  NAND2X1 U6020 ( .A(inst_data_MEM_data[154]), .B(n4966), .Y(n4961) );
  OAI21X1 U6021 ( .A(n4965), .B(n5109), .C(n4961), .Y(n2560) );
  NAND2X1 U6022 ( .A(inst_data_MEM_data[155]), .B(n4966), .Y(n4962) );
  OAI21X1 U6023 ( .A(n4965), .B(n5111), .C(n4962), .Y(n2559) );
  NAND2X1 U6024 ( .A(inst_data_MEM_data[156]), .B(n4966), .Y(n4963) );
  OAI21X1 U6025 ( .A(n4965), .B(n5114), .C(n4963), .Y(n2558) );
  NAND2X1 U6026 ( .A(inst_data_MEM_data[157]), .B(n4966), .Y(n4964) );
  OAI21X1 U6027 ( .A(n4965), .B(n5116), .C(n4964), .Y(n2557) );
  NAND2X1 U6028 ( .A(inst_data_MEM_data[158]), .B(n4966), .Y(n4967) );
  OAI21X1 U6029 ( .A(n4968), .B(n5118), .C(n4967), .Y(n2556) );
  NAND2X1 U6030 ( .A(inst_data_MEM_data[127]), .B(n4754), .Y(n4969) );
  OAI21X1 U6031 ( .A(n5067), .B(n5002), .C(n4969), .Y(n2555) );
  NAND2X1 U6032 ( .A(inst_data_MEM_data[99]), .B(n4754), .Y(n4970) );
  OAI21X1 U6033 ( .A(n4971), .B(n5002), .C(n4970), .Y(n2554) );
  NAND2X1 U6034 ( .A(inst_data_MEM_data[100]), .B(n4754), .Y(n4972) );
  OAI21X1 U6035 ( .A(n4973), .B(n5002), .C(n4972), .Y(n2553) );
  NAND2X1 U6036 ( .A(inst_data_MEM_data[101]), .B(n4754), .Y(n4974) );
  OAI21X1 U6037 ( .A(n4975), .B(n5002), .C(n4974), .Y(n2552) );
  NAND2X1 U6038 ( .A(inst_data_MEM_data[102]), .B(n4754), .Y(n4976) );
  OAI21X1 U6039 ( .A(n5069), .B(n5002), .C(n4976), .Y(n2551) );
  NAND2X1 U6040 ( .A(inst_data_MEM_data[103]), .B(n4754), .Y(n4977) );
  OAI21X1 U6041 ( .A(n5071), .B(n5002), .C(n4977), .Y(n2550) );
  NAND2X1 U6042 ( .A(inst_data_MEM_data[104]), .B(n4754), .Y(n4978) );
  OAI21X1 U6043 ( .A(n5073), .B(n5002), .C(n4978), .Y(n2549) );
  NAND2X1 U6044 ( .A(inst_data_MEM_data[105]), .B(n4754), .Y(n4979) );
  OAI21X1 U6045 ( .A(n5075), .B(n5002), .C(n4979), .Y(n2548) );
  NAND2X1 U6046 ( .A(inst_data_MEM_data[106]), .B(n4754), .Y(n4980) );
  OAI21X1 U6047 ( .A(n5077), .B(n5002), .C(n4980), .Y(n2547) );
  NAND2X1 U6048 ( .A(inst_data_MEM_data[107]), .B(n4754), .Y(n4981) );
  OAI21X1 U6049 ( .A(n5079), .B(n5002), .C(n4981), .Y(n2546) );
  NAND2X1 U6050 ( .A(inst_data_MEM_data[108]), .B(n5000), .Y(n4982) );
  OAI21X1 U6051 ( .A(n5081), .B(n5002), .C(n4982), .Y(n2545) );
  NAND2X1 U6052 ( .A(inst_data_MEM_data[109]), .B(n5000), .Y(n4983) );
  OAI21X1 U6053 ( .A(n5083), .B(n5002), .C(n4983), .Y(n2544) );
  NAND2X1 U6054 ( .A(inst_data_MEM_data[110]), .B(n4754), .Y(n4984) );
  OAI21X1 U6055 ( .A(n5085), .B(n5002), .C(n4984), .Y(n2543) );
  NAND2X1 U6056 ( .A(inst_data_MEM_data[111]), .B(n5000), .Y(n4985) );
  OAI21X1 U6057 ( .A(n5087), .B(n5002), .C(n4985), .Y(n2542) );
  NAND2X1 U6058 ( .A(inst_data_MEM_data[112]), .B(n5000), .Y(n4986) );
  OAI21X1 U6059 ( .A(n5089), .B(n5002), .C(n4986), .Y(n2541) );
  NAND2X1 U6060 ( .A(inst_data_MEM_data[113]), .B(n4754), .Y(n4987) );
  OAI21X1 U6061 ( .A(n5091), .B(n5002), .C(n4987), .Y(n2540) );
  NAND2X1 U6062 ( .A(inst_data_MEM_data[114]), .B(n4754), .Y(n4988) );
  OAI21X1 U6063 ( .A(n5093), .B(n5002), .C(n4988), .Y(n2539) );
  NAND2X1 U6064 ( .A(inst_data_MEM_data[115]), .B(n4754), .Y(n4989) );
  OAI21X1 U6065 ( .A(n5095), .B(n5002), .C(n4989), .Y(n2538) );
  NAND2X1 U6066 ( .A(inst_data_MEM_data[116]), .B(n4754), .Y(n4990) );
  OAI21X1 U6067 ( .A(n5097), .B(n5002), .C(n4990), .Y(n2537) );
  NAND2X1 U6068 ( .A(inst_data_MEM_data[117]), .B(n4754), .Y(n4991) );
  OAI21X1 U6069 ( .A(n5099), .B(n5002), .C(n4991), .Y(n2536) );
  NAND2X1 U6070 ( .A(inst_data_MEM_data[118]), .B(n4754), .Y(n4992) );
  OAI21X1 U6071 ( .A(n5101), .B(n5002), .C(n4992), .Y(n2535) );
  NAND2X1 U6072 ( .A(inst_data_MEM_data[119]), .B(n4754), .Y(n4993) );
  OAI21X1 U6073 ( .A(n5103), .B(n5002), .C(n4993), .Y(n2534) );
  NAND2X1 U6074 ( .A(inst_data_MEM_data[120]), .B(n5000), .Y(n4994) );
  OAI21X1 U6075 ( .A(n5105), .B(n5002), .C(n4994), .Y(n2533) );
  NAND2X1 U6076 ( .A(inst_data_MEM_data[121]), .B(n5000), .Y(n4995) );
  OAI21X1 U6077 ( .A(n5107), .B(n5002), .C(n4995), .Y(n2532) );
  NAND2X1 U6078 ( .A(inst_data_MEM_data[122]), .B(n5000), .Y(n4996) );
  OAI21X1 U6079 ( .A(n5109), .B(n5002), .C(n4996), .Y(n2531) );
  NAND2X1 U6080 ( .A(inst_data_MEM_data[123]), .B(n5000), .Y(n4997) );
  OAI21X1 U6081 ( .A(n5111), .B(n5002), .C(n4997), .Y(n2530) );
  NAND2X1 U6082 ( .A(inst_data_MEM_data[124]), .B(n5000), .Y(n4998) );
  OAI21X1 U6083 ( .A(n5114), .B(n5002), .C(n4998), .Y(n2529) );
  NAND2X1 U6084 ( .A(inst_data_MEM_data[125]), .B(n5000), .Y(n4999) );
  OAI21X1 U6085 ( .A(n5116), .B(n5002), .C(n4999), .Y(n2528) );
  NAND2X1 U6086 ( .A(inst_data_MEM_data[126]), .B(n5000), .Y(n5001) );
  OAI21X1 U6087 ( .A(n5118), .B(n5002), .C(n5001), .Y(n2527) );
  INVX1 U6088 ( .A(inst_data_MEM_data[253]), .Y(n5004) );
  NAND2X1 U6089 ( .A(n5062), .B(write_mem_data_MEM[29]), .Y(n5003) );
  OAI21X1 U6090 ( .A(n5065), .B(n5004), .C(n5003), .Y(n2526) );
  INVX1 U6091 ( .A(write_mem_data_MEM[0]), .Y(n5006) );
  NAND2X1 U6092 ( .A(inst_data_MEM_data[224]), .B(n5009), .Y(n5005) );
  OAI21X1 U6093 ( .A(n5006), .B(n5014), .C(n5005), .Y(n2525) );
  INVX1 U6094 ( .A(write_mem_data_MEM[1]), .Y(n5008) );
  NAND2X1 U6095 ( .A(inst_data_MEM_data[225]), .B(n5009), .Y(n5007) );
  OAI21X1 U6096 ( .A(n5008), .B(n5014), .C(n5007), .Y(n2524) );
  INVX1 U6097 ( .A(write_mem_data_MEM[2]), .Y(n5011) );
  NAND2X1 U6098 ( .A(inst_data_MEM_data[226]), .B(n5009), .Y(n5010) );
  OAI21X1 U6099 ( .A(n5011), .B(n5014), .C(n5010), .Y(n2523) );
  INVX1 U6100 ( .A(inst_data_MEM_data[228]), .Y(n5013) );
  NAND2X1 U6101 ( .A(n5062), .B(write_mem_data_MEM[4]), .Y(n5012) );
  OAI21X1 U6102 ( .A(n5065), .B(n5013), .C(n5012), .Y(n2521) );
  INVX1 U6103 ( .A(inst_data_MEM_data[229]), .Y(n5016) );
  NAND2X1 U6104 ( .A(n5062), .B(write_mem_data_MEM[5]), .Y(n5015) );
  OAI21X1 U6105 ( .A(n5065), .B(n5016), .C(n5015), .Y(n2520) );
  INVX1 U6106 ( .A(inst_data_MEM_data[230]), .Y(n5018) );
  NAND2X1 U6107 ( .A(n5062), .B(write_mem_data_MEM[6]), .Y(n5017) );
  OAI21X1 U6108 ( .A(n5065), .B(n5018), .C(n5017), .Y(n2519) );
  INVX1 U6109 ( .A(inst_data_MEM_data[231]), .Y(n5020) );
  NAND2X1 U6110 ( .A(n5062), .B(write_mem_data_MEM[7]), .Y(n5019) );
  OAI21X1 U6111 ( .A(n5065), .B(n5020), .C(n5019), .Y(n2518) );
  INVX1 U6112 ( .A(inst_data_MEM_data[232]), .Y(n5022) );
  NAND2X1 U6113 ( .A(n5062), .B(write_mem_data_MEM[8]), .Y(n5021) );
  OAI21X1 U6114 ( .A(n5065), .B(n5022), .C(n5021), .Y(n2517) );
  INVX1 U6115 ( .A(inst_data_MEM_data[233]), .Y(n5024) );
  NAND2X1 U6116 ( .A(n5062), .B(write_mem_data_MEM[9]), .Y(n5023) );
  OAI21X1 U6117 ( .A(n5065), .B(n5024), .C(n5023), .Y(n2516) );
  INVX1 U6118 ( .A(inst_data_MEM_data[234]), .Y(n5026) );
  NAND2X1 U6119 ( .A(n5062), .B(write_mem_data_MEM[10]), .Y(n5025) );
  OAI21X1 U6120 ( .A(n5065), .B(n5026), .C(n5025), .Y(n2515) );
  INVX1 U6121 ( .A(inst_data_MEM_data[235]), .Y(n5028) );
  NAND2X1 U6122 ( .A(n5062), .B(write_mem_data_MEM[11]), .Y(n5027) );
  OAI21X1 U6123 ( .A(n5065), .B(n5028), .C(n5027), .Y(n2514) );
  INVX1 U6124 ( .A(inst_data_MEM_data[236]), .Y(n5030) );
  NAND2X1 U6125 ( .A(n5062), .B(write_mem_data_MEM[12]), .Y(n5029) );
  OAI21X1 U6126 ( .A(n5065), .B(n5030), .C(n5029), .Y(n2513) );
  INVX1 U6127 ( .A(inst_data_MEM_data[237]), .Y(n5032) );
  NAND2X1 U6128 ( .A(n5062), .B(write_mem_data_MEM[13]), .Y(n5031) );
  OAI21X1 U6129 ( .A(n5065), .B(n5032), .C(n5031), .Y(n2512) );
  INVX1 U6130 ( .A(inst_data_MEM_data[238]), .Y(n5034) );
  NAND2X1 U6131 ( .A(n5062), .B(write_mem_data_MEM[14]), .Y(n5033) );
  OAI21X1 U6132 ( .A(n5065), .B(n5034), .C(n5033), .Y(n2511) );
  INVX1 U6133 ( .A(inst_data_MEM_data[239]), .Y(n5036) );
  NAND2X1 U6134 ( .A(n5062), .B(write_mem_data_MEM[15]), .Y(n5035) );
  OAI21X1 U6135 ( .A(n5065), .B(n5036), .C(n5035), .Y(n2510) );
  INVX1 U6136 ( .A(inst_data_MEM_data[240]), .Y(n5038) );
  NAND2X1 U6137 ( .A(n5062), .B(write_mem_data_MEM[16]), .Y(n5037) );
  OAI21X1 U6138 ( .A(n5065), .B(n5038), .C(n5037), .Y(n2509) );
  INVX1 U6139 ( .A(inst_data_MEM_data[241]), .Y(n5040) );
  NAND2X1 U6140 ( .A(n5062), .B(write_mem_data_MEM[17]), .Y(n5039) );
  OAI21X1 U6141 ( .A(n5061), .B(n5040), .C(n5039), .Y(n2508) );
  INVX1 U6142 ( .A(inst_data_MEM_data[242]), .Y(n5042) );
  NAND2X1 U6143 ( .A(n5062), .B(write_mem_data_MEM[18]), .Y(n5041) );
  OAI21X1 U6144 ( .A(n5061), .B(n5042), .C(n5041), .Y(n2507) );
  INVX1 U6145 ( .A(inst_data_MEM_data[243]), .Y(n5044) );
  NAND2X1 U6146 ( .A(n5062), .B(write_mem_data_MEM[19]), .Y(n5043) );
  OAI21X1 U6147 ( .A(n5061), .B(n5044), .C(n5043), .Y(n2506) );
  INVX1 U6148 ( .A(inst_data_MEM_data[244]), .Y(n5046) );
  NAND2X1 U6149 ( .A(n5062), .B(write_mem_data_MEM[20]), .Y(n5045) );
  OAI21X1 U6150 ( .A(n5061), .B(n5046), .C(n5045), .Y(n2505) );
  INVX1 U6151 ( .A(inst_data_MEM_data[245]), .Y(n5048) );
  NAND2X1 U6152 ( .A(n5062), .B(write_mem_data_MEM[21]), .Y(n5047) );
  OAI21X1 U6153 ( .A(n5061), .B(n5048), .C(n5047), .Y(n2504) );
  INVX1 U6154 ( .A(inst_data_MEM_data[246]), .Y(n5050) );
  NAND2X1 U6155 ( .A(n5062), .B(write_mem_data_MEM[22]), .Y(n5049) );
  OAI21X1 U6156 ( .A(n5061), .B(n5050), .C(n5049), .Y(n2503) );
  INVX1 U6157 ( .A(inst_data_MEM_data[247]), .Y(n5052) );
  NAND2X1 U6158 ( .A(n5062), .B(write_mem_data_MEM[23]), .Y(n5051) );
  OAI21X1 U6159 ( .A(n5061), .B(n5052), .C(n5051), .Y(n2502) );
  INVX1 U6160 ( .A(inst_data_MEM_data[248]), .Y(n5054) );
  NAND2X1 U6161 ( .A(n5062), .B(write_mem_data_MEM[24]), .Y(n5053) );
  OAI21X1 U6162 ( .A(n5061), .B(n5054), .C(n5053), .Y(n2501) );
  INVX1 U6163 ( .A(inst_data_MEM_data[249]), .Y(n5056) );
  NAND2X1 U6164 ( .A(n5062), .B(write_mem_data_MEM[25]), .Y(n5055) );
  OAI21X1 U6165 ( .A(n5061), .B(n5056), .C(n5055), .Y(n2500) );
  INVX1 U6166 ( .A(inst_data_MEM_data[250]), .Y(n5058) );
  NAND2X1 U6167 ( .A(n5062), .B(write_mem_data_MEM[26]), .Y(n5057) );
  OAI21X1 U6168 ( .A(n5061), .B(n5058), .C(n5057), .Y(n2499) );
  INVX1 U6169 ( .A(inst_data_MEM_data[251]), .Y(n5060) );
  NAND2X1 U6170 ( .A(n5062), .B(write_mem_data_MEM[27]), .Y(n5059) );
  OAI21X1 U6171 ( .A(n5061), .B(n5060), .C(n5059), .Y(n2498) );
  INVX1 U6172 ( .A(inst_data_MEM_data[252]), .Y(n5064) );
  NAND2X1 U6173 ( .A(n5062), .B(write_mem_data_MEM[28]), .Y(n5063) );
  OAI21X1 U6174 ( .A(n5065), .B(n5064), .C(n5063), .Y(n2497) );
  NAND2X1 U6175 ( .A(inst_data_MEM_data[223]), .B(n4878), .Y(n5066) );
  OAI21X1 U6176 ( .A(n5119), .B(n5067), .C(n5066), .Y(n2496) );
  NAND2X1 U6177 ( .A(inst_data_MEM_data[198]), .B(n4878), .Y(n5068) );
  OAI21X1 U6178 ( .A(n5119), .B(n5069), .C(n5068), .Y(n2495) );
  NAND2X1 U6179 ( .A(inst_data_MEM_data[199]), .B(n4878), .Y(n5070) );
  OAI21X1 U6180 ( .A(n5119), .B(n5071), .C(n5070), .Y(n2494) );
  NAND2X1 U6181 ( .A(inst_data_MEM_data[200]), .B(n4878), .Y(n5072) );
  OAI21X1 U6182 ( .A(n5119), .B(n5073), .C(n5072), .Y(n2493) );
  NAND2X1 U6183 ( .A(inst_data_MEM_data[201]), .B(n4878), .Y(n5074) );
  OAI21X1 U6184 ( .A(n5119), .B(n5075), .C(n5074), .Y(n2492) );
  NAND2X1 U6185 ( .A(inst_data_MEM_data[202]), .B(n4878), .Y(n5076) );
  OAI21X1 U6186 ( .A(n5119), .B(n5077), .C(n5076), .Y(n2491) );
  NAND2X1 U6187 ( .A(inst_data_MEM_data[203]), .B(n4878), .Y(n5078) );
  OAI21X1 U6188 ( .A(n5119), .B(n5079), .C(n5078), .Y(n2490) );
  NAND2X1 U6189 ( .A(inst_data_MEM_data[204]), .B(n4878), .Y(n5080) );
  OAI21X1 U6190 ( .A(n5119), .B(n5081), .C(n5080), .Y(n2489) );
  NAND2X1 U6191 ( .A(inst_data_MEM_data[205]), .B(n4878), .Y(n5082) );
  OAI21X1 U6192 ( .A(n5119), .B(n5083), .C(n5082), .Y(n2488) );
  NAND2X1 U6193 ( .A(inst_data_MEM_data[206]), .B(n5112), .Y(n5084) );
  OAI21X1 U6194 ( .A(n5119), .B(n5085), .C(n5084), .Y(n2487) );
  NAND2X1 U6195 ( .A(inst_data_MEM_data[207]), .B(n5112), .Y(n5086) );
  OAI21X1 U6196 ( .A(n5119), .B(n5087), .C(n5086), .Y(n2486) );
  NAND2X1 U6197 ( .A(inst_data_MEM_data[208]), .B(n5112), .Y(n5088) );
  OAI21X1 U6198 ( .A(n5119), .B(n5089), .C(n5088), .Y(n2485) );
  NAND2X1 U6199 ( .A(inst_data_MEM_data[209]), .B(n5112), .Y(n5090) );
  OAI21X1 U6200 ( .A(n5119), .B(n5091), .C(n5090), .Y(n2484) );
  NAND2X1 U6201 ( .A(inst_data_MEM_data[210]), .B(n5112), .Y(n5092) );
  OAI21X1 U6202 ( .A(n5119), .B(n5093), .C(n5092), .Y(n2483) );
  NAND2X1 U6203 ( .A(inst_data_MEM_data[211]), .B(n5112), .Y(n5094) );
  OAI21X1 U6204 ( .A(n5119), .B(n5095), .C(n5094), .Y(n2482) );
  NAND2X1 U6205 ( .A(inst_data_MEM_data[212]), .B(n5112), .Y(n5096) );
  OAI21X1 U6206 ( .A(n5119), .B(n5097), .C(n5096), .Y(n2481) );
  NAND2X1 U6207 ( .A(inst_data_MEM_data[213]), .B(n5112), .Y(n5098) );
  OAI21X1 U6208 ( .A(n5119), .B(n5099), .C(n5098), .Y(n2480) );
  NAND2X1 U6209 ( .A(inst_data_MEM_data[214]), .B(n5112), .Y(n5100) );
  OAI21X1 U6210 ( .A(n5119), .B(n5101), .C(n5100), .Y(n2479) );
  NAND2X1 U6211 ( .A(inst_data_MEM_data[215]), .B(n4878), .Y(n5102) );
  OAI21X1 U6212 ( .A(n5119), .B(n5103), .C(n5102), .Y(n2478) );
  NAND2X1 U6213 ( .A(inst_data_MEM_data[216]), .B(n5112), .Y(n5104) );
  OAI21X1 U6214 ( .A(n5119), .B(n5105), .C(n5104), .Y(n2477) );
  NAND2X1 U6215 ( .A(inst_data_MEM_data[217]), .B(n4878), .Y(n5106) );
  OAI21X1 U6216 ( .A(n5119), .B(n5107), .C(n5106), .Y(n2476) );
  NAND2X1 U6217 ( .A(inst_data_MEM_data[218]), .B(n4878), .Y(n5108) );
  OAI21X1 U6218 ( .A(n5119), .B(n5109), .C(n5108), .Y(n2475) );
  NAND2X1 U6219 ( .A(inst_data_MEM_data[219]), .B(n5112), .Y(n5110) );
  OAI21X1 U6220 ( .A(n5119), .B(n5111), .C(n5110), .Y(n2474) );
  NAND2X1 U6221 ( .A(inst_data_MEM_data[220]), .B(n5112), .Y(n5113) );
  OAI21X1 U6222 ( .A(n5119), .B(n5114), .C(n5113), .Y(n2473) );
  NAND2X1 U6223 ( .A(inst_data_MEM_data[221]), .B(n4878), .Y(n5115) );
  OAI21X1 U6224 ( .A(n5119), .B(n5116), .C(n5115), .Y(n2472) );
  NAND2X1 U6225 ( .A(inst_data_MEM_data[222]), .B(n4878), .Y(n5117) );
  OAI21X1 U6226 ( .A(n5119), .B(n5118), .C(n5117), .Y(n2471) );
  INVX1 U6227 ( .A(inst_register_registers[253]), .Y(n5123) );
  NAND2X1 U6228 ( .A(n5202), .B(reg_write_address_WB[0]), .Y(n5243) );
  NOR2X1 U6229 ( .A(n5428), .B(n5243), .Y(n5315) );
  NAND2X1 U6230 ( .A(reg_write_address_WB[2]), .B(n5315), .Y(n5234) );
  AND2X2 U6231 ( .A(n3066), .B(n5120), .Y(n5155) );
  NAND2X1 U6232 ( .A(n3066), .B(n5122), .Y(n5493) );
  OAI22X1 U6233 ( .A(n5123), .B(n2811), .C(n5493), .D(n5120), .Y(n2470) );
  INVX1 U6234 ( .A(inst_register_registers[224]), .Y(n5125) );
  NAND2X1 U6235 ( .A(n2815), .B(n5124), .Y(n5433) );
  OAI22X1 U6236 ( .A(n5125), .B(n2811), .C(n5120), .D(n5433), .Y(n2469) );
  INVX1 U6237 ( .A(inst_register_registers[225]), .Y(n5128) );
  NAND2X1 U6238 ( .A(n2815), .B(n5127), .Y(n5435) );
  OAI22X1 U6239 ( .A(n5128), .B(n2811), .C(n5120), .D(n5435), .Y(n2468) );
  INVX1 U6240 ( .A(inst_register_registers[226]), .Y(n5131) );
  INVX1 U6241 ( .A(n5129), .Y(n5130) );
  NAND2X1 U6242 ( .A(n2815), .B(n5130), .Y(n5438) );
  OAI22X1 U6243 ( .A(n5131), .B(n2811), .C(n5120), .D(n5438), .Y(n2467) );
  INVX1 U6244 ( .A(inst_register_registers[227]), .Y(n5134) );
  INVX1 U6245 ( .A(n5132), .Y(n5133) );
  NAND2X1 U6246 ( .A(n2815), .B(n5133), .Y(n5440) );
  OAI22X1 U6247 ( .A(n5134), .B(n2811), .C(n5120), .D(n5440), .Y(n2466) );
  INVX1 U6248 ( .A(inst_register_registers[228]), .Y(n5137) );
  NAND2X1 U6249 ( .A(n2815), .B(n5136), .Y(n5442) );
  OAI22X1 U6250 ( .A(n5137), .B(n2811), .C(n5120), .D(n5442), .Y(n2465) );
  INVX1 U6251 ( .A(inst_register_registers[229]), .Y(n5140) );
  INVX1 U6252 ( .A(n5138), .Y(n5139) );
  NAND2X1 U6253 ( .A(n3066), .B(n5139), .Y(n5444) );
  OAI22X1 U6254 ( .A(n5140), .B(n2811), .C(n5120), .D(n5444), .Y(n2464) );
  INVX1 U6255 ( .A(inst_register_registers[230]), .Y(n5143) );
  INVX1 U6256 ( .A(n5141), .Y(n5142) );
  NAND2X1 U6257 ( .A(n3066), .B(n5142), .Y(n5446) );
  OAI22X1 U6258 ( .A(n5143), .B(n2811), .C(n5234), .D(n5446), .Y(n2463) );
  INVX1 U6259 ( .A(inst_register_registers[231]), .Y(n5146) );
  NAND2X1 U6260 ( .A(n2815), .B(n5145), .Y(n5448) );
  OAI22X1 U6261 ( .A(n5146), .B(n2811), .C(n5234), .D(n5448), .Y(n2462) );
  INVX1 U6262 ( .A(inst_register_registers[232]), .Y(n5148) );
  NAND2X1 U6263 ( .A(n2815), .B(n5147), .Y(n5450) );
  OAI22X1 U6264 ( .A(n5148), .B(n2811), .C(n5234), .D(n5450), .Y(n2461) );
  INVX1 U6265 ( .A(inst_register_registers[233]), .Y(n5151) );
  NAND2X1 U6266 ( .A(n2815), .B(n5150), .Y(n5452) );
  OAI22X1 U6267 ( .A(n5151), .B(n2811), .C(n5234), .D(n5452), .Y(n2460) );
  INVX1 U6268 ( .A(inst_register_registers[234]), .Y(n5154) );
  INVX1 U6269 ( .A(n5152), .Y(n5153) );
  NAND2X1 U6270 ( .A(n2815), .B(n5153), .Y(n5454) );
  OAI22X1 U6271 ( .A(n5154), .B(n2811), .C(n5234), .D(n5454), .Y(n2459) );
  INVX1 U6272 ( .A(inst_register_registers[235]), .Y(n5158) );
  INVX1 U6273 ( .A(n5156), .Y(n5157) );
  NAND2X1 U6274 ( .A(n3066), .B(n5157), .Y(n5456) );
  OAI22X1 U6275 ( .A(n5158), .B(n2811), .C(n5234), .D(n5456), .Y(n2458) );
  INVX1 U6276 ( .A(inst_register_registers[236]), .Y(n5161) );
  INVX1 U6277 ( .A(n5159), .Y(n5160) );
  NAND2X1 U6278 ( .A(n2815), .B(n5160), .Y(n5458) );
  OAI22X1 U6279 ( .A(n5161), .B(n2811), .C(n5120), .D(n5458), .Y(n2457) );
  INVX1 U6280 ( .A(inst_register_registers[237]), .Y(n5164) );
  NAND2X1 U6281 ( .A(n2815), .B(n5163), .Y(n5460) );
  OAI22X1 U6282 ( .A(n5164), .B(n2811), .C(n5120), .D(n5460), .Y(n2456) );
  INVX1 U6283 ( .A(inst_register_registers[238]), .Y(n5166) );
  NAND2X1 U6284 ( .A(n2815), .B(n5165), .Y(n5462) );
  OAI22X1 U6285 ( .A(n5166), .B(n2811), .C(n5120), .D(n5462), .Y(n2455) );
  INVX1 U6286 ( .A(inst_register_registers[239]), .Y(n5168) );
  NAND2X1 U6287 ( .A(n2815), .B(n5167), .Y(n5464) );
  OAI22X1 U6288 ( .A(n5168), .B(n2811), .C(n5120), .D(n5464), .Y(n2454) );
  INVX1 U6289 ( .A(inst_register_registers[240]), .Y(n5170) );
  NAND2X1 U6290 ( .A(n2815), .B(n5169), .Y(n5466) );
  OAI22X1 U6291 ( .A(n5170), .B(n2811), .C(n5234), .D(n5466), .Y(n2453) );
  INVX1 U6292 ( .A(inst_register_registers[241]), .Y(n5173) );
  NAND2X1 U6293 ( .A(n2815), .B(n5172), .Y(n5468) );
  OAI22X1 U6294 ( .A(n5173), .B(n2811), .C(n5120), .D(n5468), .Y(n2452) );
  INVX1 U6295 ( .A(inst_register_registers[242]), .Y(n5175) );
  NAND2X1 U6296 ( .A(n2815), .B(n5174), .Y(n5470) );
  OAI22X1 U6297 ( .A(n5175), .B(n2811), .C(n5120), .D(n5470), .Y(n2451) );
  INVX1 U6298 ( .A(inst_register_registers[243]), .Y(n5177) );
  NAND2X1 U6299 ( .A(n2815), .B(n5176), .Y(n5472) );
  OAI22X1 U6300 ( .A(n5177), .B(n2811), .C(n5120), .D(n5472), .Y(n2450) );
  INVX1 U6301 ( .A(inst_register_registers[244]), .Y(n5179) );
  NAND2X1 U6302 ( .A(n2815), .B(n5178), .Y(n5474) );
  OAI22X1 U6303 ( .A(n5179), .B(n2811), .C(n5120), .D(n5474), .Y(n2449) );
  INVX1 U6304 ( .A(inst_register_registers[245]), .Y(n5181) );
  NAND2X1 U6305 ( .A(n2815), .B(n5180), .Y(n5476) );
  OAI22X1 U6306 ( .A(n5181), .B(n2811), .C(n5120), .D(n5476), .Y(n2448) );
  INVX1 U6307 ( .A(inst_register_registers[246]), .Y(n5183) );
  NAND2X1 U6308 ( .A(n2815), .B(n5182), .Y(n5478) );
  OAI22X1 U6309 ( .A(n5183), .B(n2811), .C(n5120), .D(n5478), .Y(n2447) );
  INVX1 U6310 ( .A(inst_register_registers[247]), .Y(n5185) );
  NAND2X1 U6311 ( .A(n2815), .B(n5184), .Y(n5480) );
  OAI22X1 U6312 ( .A(n5185), .B(n2811), .C(n5234), .D(n5480), .Y(n2446) );
  INVX1 U6313 ( .A(inst_register_registers[248]), .Y(n5188) );
  INVX1 U6314 ( .A(n5186), .Y(n5187) );
  NAND2X1 U6315 ( .A(n3066), .B(n5187), .Y(n5482) );
  OAI22X1 U6316 ( .A(n5188), .B(n2811), .C(n5234), .D(n5482), .Y(n2445) );
  INVX1 U6317 ( .A(inst_register_registers[249]), .Y(n5191) );
  NAND2X1 U6318 ( .A(n3066), .B(n5190), .Y(n5484) );
  OAI22X1 U6319 ( .A(n5191), .B(n2811), .C(n5234), .D(n5484), .Y(n2444) );
  INVX1 U6320 ( .A(inst_register_registers[250]), .Y(n5194) );
  NAND2X1 U6321 ( .A(n3066), .B(n5193), .Y(n5487) );
  OAI22X1 U6322 ( .A(n5194), .B(n2811), .C(n5234), .D(n5487), .Y(n2443) );
  INVX1 U6323 ( .A(inst_register_registers[251]), .Y(n5197) );
  NAND2X1 U6324 ( .A(n3066), .B(n5196), .Y(n5489) );
  OAI22X1 U6325 ( .A(n5197), .B(n2811), .C(n5120), .D(n5489), .Y(n2442) );
  INVX1 U6326 ( .A(inst_register_registers[252]), .Y(n5200) );
  NAND2X1 U6327 ( .A(n3066), .B(n5199), .Y(n5491) );
  OAI22X1 U6328 ( .A(n5200), .B(n2811), .C(n5120), .D(n5491), .Y(n2441) );
  INVX1 U6329 ( .A(inst_register_registers[223]), .Y(n5205) );
  NAND2X1 U6330 ( .A(n5202), .B(n5201), .Y(n5353) );
  NOR2X1 U6331 ( .A(n5391), .B(n5353), .Y(n5279) );
  NAND2X1 U6332 ( .A(reg_write_address_WB[1]), .B(n5279), .Y(n5240) );
  AND2X2 U6333 ( .A(n3066), .B(n5203), .Y(n5209) );
  NAND2X1 U6334 ( .A(n2815), .B(n5204), .Y(n5431) );
  OAI22X1 U6335 ( .A(n5205), .B(n2810), .C(n5431), .D(n5203), .Y(n2440) );
  INVX1 U6336 ( .A(inst_register_registers[198]), .Y(n5206) );
  OAI22X1 U6337 ( .A(n5206), .B(n2810), .C(n5446), .D(n5203), .Y(n2439) );
  INVX1 U6338 ( .A(inst_register_registers[199]), .Y(n5207) );
  OAI22X1 U6339 ( .A(n5207), .B(n2810), .C(n5448), .D(n5240), .Y(n2438) );
  INVX1 U6340 ( .A(inst_register_registers[200]), .Y(n5208) );
  OAI22X1 U6341 ( .A(n5208), .B(n2810), .C(n5450), .D(n5203), .Y(n2437) );
  INVX1 U6342 ( .A(inst_register_registers[201]), .Y(n5210) );
  OAI22X1 U6343 ( .A(n5210), .B(n2810), .C(n5452), .D(n5203), .Y(n2436) );
  INVX1 U6344 ( .A(inst_register_registers[202]), .Y(n5211) );
  OAI22X1 U6345 ( .A(n5211), .B(n2810), .C(n5454), .D(n5240), .Y(n2435) );
  INVX1 U6346 ( .A(inst_register_registers[203]), .Y(n5212) );
  OAI22X1 U6347 ( .A(n5212), .B(n2810), .C(n5456), .D(n5240), .Y(n2434) );
  INVX1 U6348 ( .A(inst_register_registers[204]), .Y(n5213) );
  OAI22X1 U6349 ( .A(n5213), .B(n2810), .C(n5458), .D(n5240), .Y(n2433) );
  INVX1 U6350 ( .A(inst_register_registers[205]), .Y(n5214) );
  OAI22X1 U6351 ( .A(n5214), .B(n2810), .C(n5460), .D(n5240), .Y(n2432) );
  INVX1 U6352 ( .A(inst_register_registers[206]), .Y(n5215) );
  OAI22X1 U6353 ( .A(n5215), .B(n2810), .C(n5462), .D(n5240), .Y(n2431) );
  INVX1 U6354 ( .A(inst_register_registers[207]), .Y(n5216) );
  OAI22X1 U6355 ( .A(n5216), .B(n2810), .C(n5464), .D(n5203), .Y(n2430) );
  INVX1 U6356 ( .A(inst_register_registers[208]), .Y(n5217) );
  OAI22X1 U6357 ( .A(n5217), .B(n2810), .C(n5466), .D(n5240), .Y(n2429) );
  INVX1 U6358 ( .A(inst_register_registers[209]), .Y(n5218) );
  OAI22X1 U6359 ( .A(n5218), .B(n2810), .C(n5468), .D(n5203), .Y(n2428) );
  INVX1 U6360 ( .A(inst_register_registers[210]), .Y(n5219) );
  OAI22X1 U6361 ( .A(n5219), .B(n2810), .C(n5470), .D(n5203), .Y(n2427) );
  INVX1 U6362 ( .A(inst_register_registers[211]), .Y(n5220) );
  OAI22X1 U6363 ( .A(n5220), .B(n2810), .C(n5472), .D(n5240), .Y(n2426) );
  INVX1 U6364 ( .A(inst_register_registers[212]), .Y(n5221) );
  OAI22X1 U6365 ( .A(n5221), .B(n2810), .C(n5474), .D(n5203), .Y(n2425) );
  INVX1 U6366 ( .A(inst_register_registers[213]), .Y(n5222) );
  OAI22X1 U6367 ( .A(n5222), .B(n2810), .C(n5476), .D(n5203), .Y(n2424) );
  INVX1 U6368 ( .A(inst_register_registers[214]), .Y(n5223) );
  OAI22X1 U6369 ( .A(n5223), .B(n2810), .C(n5478), .D(n5203), .Y(n2423) );
  INVX1 U6370 ( .A(inst_register_registers[215]), .Y(n5224) );
  AOI22X1 U6371 ( .A(n5224), .B(n5203), .C(n5480), .D(n2810), .Y(n2422) );
  INVX1 U6372 ( .A(inst_register_registers[216]), .Y(n5225) );
  AOI22X1 U6373 ( .A(n5225), .B(n5203), .C(n5482), .D(n2810), .Y(n2421) );
  INVX1 U6374 ( .A(inst_register_registers[217]), .Y(n5226) );
  OAI22X1 U6375 ( .A(n5226), .B(n2810), .C(n5484), .D(n5203), .Y(n2420) );
  INVX1 U6376 ( .A(inst_register_registers[218]), .Y(n5227) );
  AOI22X1 U6377 ( .A(n5227), .B(n5203), .C(n5487), .D(n2810), .Y(n2419) );
  INVX1 U6378 ( .A(inst_register_registers[219]), .Y(n5228) );
  OAI22X1 U6379 ( .A(n5228), .B(n2810), .C(n5489), .D(n5203), .Y(n2418) );
  INVX1 U6380 ( .A(inst_register_registers[220]), .Y(n5229) );
  OAI22X1 U6381 ( .A(n5229), .B(n2810), .C(n5491), .D(n5203), .Y(n2417) );
  INVX1 U6382 ( .A(inst_register_registers[221]), .Y(n5230) );
  OAI22X1 U6383 ( .A(n5230), .B(n2810), .C(n5493), .D(n5203), .Y(n2416) );
  INVX1 U6384 ( .A(inst_register_registers[222]), .Y(n5233) );
  NAND2X1 U6385 ( .A(n3066), .B(n5232), .Y(n5495) );
  OAI22X1 U6386 ( .A(n5233), .B(n2810), .C(n5203), .D(n5495), .Y(n2415) );
  INVX1 U6387 ( .A(inst_register_registers[254]), .Y(n5235) );
  OAI22X1 U6388 ( .A(n5235), .B(n2811), .C(n5234), .D(n5495), .Y(n2414) );
  INVX1 U6389 ( .A(inst_register_registers[197]), .Y(n5236) );
  OAI22X1 U6390 ( .A(n5236), .B(n2810), .C(n5444), .D(n5203), .Y(n2413) );
  INVX1 U6391 ( .A(inst_register_registers[192]), .Y(n5237) );
  OAI22X1 U6392 ( .A(n5237), .B(n2810), .C(n5433), .D(n5240), .Y(n2412) );
  INVX1 U6393 ( .A(inst_register_registers[193]), .Y(n5238) );
  OAI22X1 U6394 ( .A(n5238), .B(n2810), .C(n5435), .D(n5240), .Y(n2411) );
  INVX1 U6395 ( .A(inst_register_registers[194]), .Y(n5239) );
  OAI22X1 U6396 ( .A(n5239), .B(n2810), .C(n5438), .D(n5240), .Y(n2410) );
  INVX1 U6397 ( .A(inst_register_registers[195]), .Y(n5241) );
  OAI22X1 U6398 ( .A(n5241), .B(n2810), .C(n5440), .D(n5240), .Y(n2409) );
  INVX1 U6399 ( .A(inst_register_registers[196]), .Y(n5242) );
  OAI22X1 U6400 ( .A(n5242), .B(n2810), .C(n5442), .D(n5203), .Y(n2408) );
  OAI21X1 U6401 ( .A(reg_write_address_WB[1]), .B(n5243), .C(n2815), .Y(n5390)
         );
  OAI21X1 U6402 ( .A(reg_write_address_WB[2]), .B(n5392), .C(n5390), .Y(n5244)
         );
  INVX1 U6403 ( .A(inst_register_registers[191]), .Y(n5245) );
  INVX2 U6404 ( .A(n5278), .Y(n5270) );
  AOI22X1 U6405 ( .A(n5278), .B(n5431), .C(n5245), .D(n5270), .Y(n2407) );
  INVX1 U6406 ( .A(inst_register_registers[160]), .Y(n5246) );
  AOI22X1 U6407 ( .A(n5278), .B(n5433), .C(n5246), .D(n5270), .Y(n2406) );
  INVX1 U6408 ( .A(inst_register_registers[161]), .Y(n5247) );
  AOI22X1 U6409 ( .A(n5278), .B(n5435), .C(n5247), .D(n5270), .Y(n2405) );
  INVX1 U6410 ( .A(inst_register_registers[162]), .Y(n5248) );
  AOI22X1 U6411 ( .A(n5278), .B(n5438), .C(n5248), .D(n5270), .Y(n2404) );
  INVX1 U6412 ( .A(inst_register_registers[163]), .Y(n5249) );
  AOI22X1 U6413 ( .A(n5278), .B(n5440), .C(n5249), .D(n5270), .Y(n2403) );
  INVX1 U6414 ( .A(inst_register_registers[164]), .Y(n5250) );
  AOI22X1 U6415 ( .A(n5278), .B(n5442), .C(n5250), .D(n5270), .Y(n2402) );
  INVX1 U6416 ( .A(inst_register_registers[165]), .Y(n5251) );
  AOI22X1 U6417 ( .A(n5278), .B(n5444), .C(n5251), .D(n5270), .Y(n2401) );
  INVX1 U6418 ( .A(inst_register_registers[166]), .Y(n5252) );
  AOI22X1 U6419 ( .A(n5278), .B(n5446), .C(n5252), .D(n5270), .Y(n2400) );
  INVX1 U6420 ( .A(inst_register_registers[167]), .Y(n5253) );
  AOI22X1 U6421 ( .A(n5278), .B(n5448), .C(n5253), .D(n5270), .Y(n2399) );
  INVX1 U6422 ( .A(inst_register_registers[168]), .Y(n5254) );
  AOI22X1 U6423 ( .A(n5278), .B(n5450), .C(n5254), .D(n5270), .Y(n2398) );
  INVX1 U6424 ( .A(inst_register_registers[169]), .Y(n5255) );
  AOI22X1 U6425 ( .A(n5278), .B(n5452), .C(n5255), .D(n5270), .Y(n2397) );
  INVX1 U6426 ( .A(inst_register_registers[170]), .Y(n5256) );
  AOI22X1 U6427 ( .A(n5278), .B(n5454), .C(n5256), .D(n5270), .Y(n2396) );
  INVX1 U6428 ( .A(inst_register_registers[171]), .Y(n5257) );
  AOI22X1 U6429 ( .A(n5278), .B(n5456), .C(n5257), .D(n5270), .Y(n2395) );
  INVX1 U6430 ( .A(inst_register_registers[172]), .Y(n5258) );
  AOI22X1 U6431 ( .A(n5278), .B(n5458), .C(n5258), .D(n5270), .Y(n2394) );
  INVX1 U6432 ( .A(inst_register_registers[173]), .Y(n5259) );
  AOI22X1 U6433 ( .A(n5278), .B(n5460), .C(n5259), .D(n5270), .Y(n2393) );
  INVX1 U6434 ( .A(inst_register_registers[174]), .Y(n5260) );
  AOI22X1 U6435 ( .A(n5278), .B(n5462), .C(n5260), .D(n5270), .Y(n2392) );
  INVX1 U6436 ( .A(inst_register_registers[175]), .Y(n5261) );
  AOI22X1 U6437 ( .A(n5278), .B(n5464), .C(n5261), .D(n5270), .Y(n2391) );
  INVX1 U6438 ( .A(inst_register_registers[176]), .Y(n5262) );
  AOI22X1 U6439 ( .A(n5278), .B(n5466), .C(n5262), .D(n5270), .Y(n2390) );
  INVX1 U6440 ( .A(inst_register_registers[177]), .Y(n5263) );
  AOI22X1 U6441 ( .A(n5278), .B(n5468), .C(n5263), .D(n5270), .Y(n2389) );
  INVX1 U6442 ( .A(inst_register_registers[178]), .Y(n5264) );
  AOI22X1 U6443 ( .A(n5278), .B(n5470), .C(n5264), .D(n5270), .Y(n2388) );
  INVX1 U6444 ( .A(inst_register_registers[179]), .Y(n5265) );
  AOI22X1 U6445 ( .A(n5278), .B(n5472), .C(n5265), .D(n5270), .Y(n2387) );
  INVX1 U6446 ( .A(inst_register_registers[180]), .Y(n5266) );
  AOI22X1 U6447 ( .A(n5278), .B(n5474), .C(n5266), .D(n5270), .Y(n2386) );
  INVX1 U6448 ( .A(inst_register_registers[181]), .Y(n5267) );
  AOI22X1 U6449 ( .A(n5278), .B(n5476), .C(n5267), .D(n5270), .Y(n2385) );
  INVX1 U6450 ( .A(inst_register_registers[182]), .Y(n5268) );
  AOI22X1 U6451 ( .A(n5278), .B(n5478), .C(n5268), .D(n5270), .Y(n2384) );
  INVX1 U6452 ( .A(inst_register_registers[183]), .Y(n5269) );
  AOI22X1 U6453 ( .A(n5278), .B(n5480), .C(n5269), .D(n5270), .Y(n2383) );
  INVX1 U6454 ( .A(inst_register_registers[184]), .Y(n5271) );
  AOI22X1 U6455 ( .A(n5278), .B(n5482), .C(n5271), .D(n5270), .Y(n2382) );
  INVX1 U6456 ( .A(inst_register_registers[185]), .Y(n5272) );
  AOI22X1 U6457 ( .A(n5278), .B(n5484), .C(n5272), .D(n5244), .Y(n2381) );
  INVX1 U6458 ( .A(inst_register_registers[186]), .Y(n5273) );
  AOI22X1 U6459 ( .A(n5278), .B(n5487), .C(n5273), .D(n5244), .Y(n2380) );
  INVX1 U6460 ( .A(inst_register_registers[187]), .Y(n5274) );
  AOI22X1 U6461 ( .A(n5278), .B(n5489), .C(n5274), .D(n5244), .Y(n2379) );
  INVX1 U6462 ( .A(inst_register_registers[188]), .Y(n5275) );
  AOI22X1 U6463 ( .A(n5278), .B(n5491), .C(n5275), .D(n5244), .Y(n2378) );
  INVX1 U6464 ( .A(inst_register_registers[189]), .Y(n5276) );
  AOI22X1 U6465 ( .A(n5278), .B(n5493), .C(n5276), .D(n5270), .Y(n2377) );
  INVX1 U6466 ( .A(inst_register_registers[190]), .Y(n5277) );
  AOI22X1 U6467 ( .A(n5278), .B(n5495), .C(n5277), .D(n5244), .Y(n2376) );
  INVX1 U6468 ( .A(inst_register_registers[159]), .Y(n5281) );
  NAND2X1 U6469 ( .A(n5279), .B(n5428), .Y(n5313) );
  AND2X2 U6470 ( .A(n3066), .B(n5280), .Y(n5282) );
  AOI22X1 U6471 ( .A(n5281), .B(n5280), .C(n5431), .D(n2812), .Y(n2375) );
  INVX1 U6472 ( .A(inst_register_registers[128]), .Y(n5283) );
  AOI22X1 U6473 ( .A(n5283), .B(n5280), .C(n5433), .D(n2812), .Y(n2374) );
  INVX1 U6474 ( .A(inst_register_registers[129]), .Y(n5284) );
  AOI22X1 U6475 ( .A(n5284), .B(n5280), .C(n5435), .D(n2812), .Y(n2373) );
  INVX1 U6476 ( .A(inst_register_registers[130]), .Y(n5285) );
  AOI22X1 U6477 ( .A(n5285), .B(n5280), .C(n5438), .D(n2812), .Y(n2372) );
  INVX1 U6478 ( .A(inst_register_registers[131]), .Y(n5286) );
  AOI22X1 U6479 ( .A(n5286), .B(n5280), .C(n5440), .D(n2812), .Y(n2371) );
  INVX1 U6480 ( .A(inst_register_registers[132]), .Y(n5287) );
  AOI22X1 U6481 ( .A(n5287), .B(n5280), .C(n5442), .D(n2812), .Y(n2370) );
  INVX1 U6482 ( .A(inst_register_registers[133]), .Y(n5288) );
  OAI22X1 U6483 ( .A(n5288), .B(n2812), .C(n5444), .D(n5280), .Y(n2369) );
  INVX1 U6484 ( .A(inst_register_registers[134]), .Y(n5289) );
  OAI22X1 U6485 ( .A(n5289), .B(n2812), .C(n5446), .D(n5280), .Y(n2368) );
  INVX1 U6486 ( .A(inst_register_registers[135]), .Y(n5290) );
  AOI22X1 U6487 ( .A(n5290), .B(n5280), .C(n5448), .D(n2812), .Y(n2367) );
  INVX1 U6488 ( .A(inst_register_registers[136]), .Y(n5291) );
  AOI22X1 U6489 ( .A(n5291), .B(n5313), .C(n5450), .D(n2812), .Y(n2366) );
  INVX1 U6490 ( .A(inst_register_registers[137]), .Y(n5292) );
  AOI22X1 U6491 ( .A(n5292), .B(n5313), .C(n5452), .D(n2812), .Y(n2365) );
  INVX1 U6492 ( .A(inst_register_registers[138]), .Y(n5293) );
  AOI22X1 U6493 ( .A(n5293), .B(n5313), .C(n5454), .D(n2812), .Y(n2364) );
  INVX1 U6494 ( .A(inst_register_registers[139]), .Y(n5294) );
  AOI22X1 U6495 ( .A(n5294), .B(n5313), .C(n5456), .D(n2812), .Y(n2363) );
  INVX1 U6496 ( .A(inst_register_registers[140]), .Y(n5295) );
  AOI22X1 U6497 ( .A(n5295), .B(n5313), .C(n5458), .D(n2812), .Y(n2362) );
  INVX1 U6498 ( .A(inst_register_registers[141]), .Y(n5296) );
  AOI22X1 U6499 ( .A(n5296), .B(n5313), .C(n5460), .D(n2812), .Y(n2361) );
  INVX1 U6500 ( .A(inst_register_registers[142]), .Y(n5297) );
  AOI22X1 U6501 ( .A(n5297), .B(n5280), .C(n5462), .D(n2812), .Y(n2360) );
  INVX1 U6502 ( .A(inst_register_registers[143]), .Y(n5298) );
  AOI22X1 U6503 ( .A(n5298), .B(n5280), .C(n5464), .D(n2812), .Y(n2359) );
  INVX1 U6504 ( .A(inst_register_registers[144]), .Y(n5299) );
  OAI22X1 U6505 ( .A(n5299), .B(n2812), .C(n5466), .D(n5280), .Y(n2358) );
  INVX1 U6506 ( .A(inst_register_registers[145]), .Y(n5300) );
  AOI22X1 U6507 ( .A(n5300), .B(n5280), .C(n5468), .D(n2812), .Y(n2357) );
  INVX1 U6508 ( .A(inst_register_registers[146]), .Y(n5301) );
  AOI22X1 U6509 ( .A(n5301), .B(n5280), .C(n5470), .D(n2812), .Y(n2356) );
  INVX1 U6510 ( .A(inst_register_registers[147]), .Y(n5302) );
  OAI22X1 U6511 ( .A(n5302), .B(n2812), .C(n5472), .D(n5280), .Y(n2355) );
  INVX1 U6512 ( .A(inst_register_registers[148]), .Y(n5303) );
  AOI22X1 U6513 ( .A(n5303), .B(n5280), .C(n5474), .D(n2812), .Y(n2354) );
  INVX1 U6514 ( .A(inst_register_registers[149]), .Y(n5304) );
  OAI22X1 U6515 ( .A(n5304), .B(n2812), .C(n5476), .D(n5280), .Y(n2353) );
  INVX1 U6516 ( .A(inst_register_registers[150]), .Y(n5305) );
  AOI22X1 U6517 ( .A(n5305), .B(n5280), .C(n5478), .D(n2812), .Y(n2352) );
  INVX1 U6518 ( .A(inst_register_registers[151]), .Y(n5306) );
  OAI22X1 U6519 ( .A(n5306), .B(n2812), .C(n5480), .D(n5313), .Y(n2351) );
  INVX1 U6520 ( .A(inst_register_registers[152]), .Y(n5307) );
  AOI22X1 U6521 ( .A(n5307), .B(n5313), .C(n5482), .D(n2812), .Y(n2350) );
  INVX1 U6522 ( .A(inst_register_registers[153]), .Y(n5308) );
  AOI22X1 U6523 ( .A(n5308), .B(n5313), .C(n5484), .D(n2812), .Y(n2349) );
  INVX1 U6524 ( .A(inst_register_registers[154]), .Y(n5309) );
  OAI22X1 U6525 ( .A(n5309), .B(n2812), .C(n5487), .D(n5313), .Y(n2348) );
  INVX1 U6526 ( .A(inst_register_registers[155]), .Y(n5310) );
  OAI22X1 U6527 ( .A(n5310), .B(n2812), .C(n5489), .D(n5280), .Y(n2347) );
  INVX1 U6528 ( .A(inst_register_registers[156]), .Y(n5311) );
  OAI22X1 U6529 ( .A(n5311), .B(n2812), .C(n5491), .D(n5313), .Y(n2346) );
  INVX1 U6530 ( .A(inst_register_registers[157]), .Y(n5312) );
  OAI22X1 U6531 ( .A(n5312), .B(n2812), .C(n5493), .D(n5280), .Y(n2345) );
  INVX1 U6532 ( .A(inst_register_registers[158]), .Y(n5314) );
  OAI22X1 U6533 ( .A(n5314), .B(n2812), .C(n5495), .D(n5313), .Y(n2344) );
  INVX1 U6534 ( .A(inst_register_registers[127]), .Y(n5318) );
  NAND2X1 U6535 ( .A(n5315), .B(n5391), .Y(n5351) );
  NAND2X1 U6536 ( .A(n2815), .B(n5316), .Y(n5345) );
  OAI22X1 U6537 ( .A(n5318), .B(n5317), .C(n5431), .D(n5316), .Y(n2343) );
  INVX1 U6538 ( .A(inst_register_registers[99]), .Y(n5319) );
  OAI22X1 U6539 ( .A(n5319), .B(n5317), .C(n5440), .D(n5316), .Y(n2342) );
  INVX1 U6540 ( .A(inst_register_registers[100]), .Y(n5320) );
  OAI22X1 U6541 ( .A(n5320), .B(n5317), .C(n5442), .D(n5316), .Y(n2341) );
  INVX1 U6542 ( .A(inst_register_registers[101]), .Y(n5321) );
  OAI22X1 U6543 ( .A(n5321), .B(n5317), .C(n5444), .D(n5316), .Y(n2340) );
  INVX1 U6544 ( .A(inst_register_registers[102]), .Y(n5322) );
  OAI22X1 U6545 ( .A(n5322), .B(n5317), .C(n5446), .D(n5316), .Y(n2339) );
  INVX1 U6546 ( .A(inst_register_registers[103]), .Y(n5323) );
  OAI22X1 U6547 ( .A(n5323), .B(n5317), .C(n5448), .D(n5316), .Y(n2338) );
  INVX1 U6548 ( .A(inst_register_registers[104]), .Y(n5324) );
  OAI22X1 U6549 ( .A(n5324), .B(n5317), .C(n5450), .D(n5316), .Y(n2337) );
  INVX1 U6550 ( .A(inst_register_registers[105]), .Y(n5325) );
  OAI22X1 U6551 ( .A(n5325), .B(n5317), .C(n5452), .D(n5316), .Y(n2336) );
  INVX1 U6552 ( .A(inst_register_registers[106]), .Y(n5326) );
  OAI22X1 U6553 ( .A(n5326), .B(n5317), .C(n5454), .D(n5351), .Y(n2335) );
  INVX1 U6554 ( .A(inst_register_registers[107]), .Y(n5327) );
  OAI22X1 U6555 ( .A(n5327), .B(n5317), .C(n5456), .D(n5351), .Y(n2334) );
  INVX1 U6556 ( .A(inst_register_registers[108]), .Y(n5328) );
  OAI22X1 U6557 ( .A(n5328), .B(n5317), .C(n5458), .D(n5351), .Y(n2333) );
  INVX1 U6558 ( .A(inst_register_registers[109]), .Y(n5329) );
  OAI22X1 U6559 ( .A(n5329), .B(n5317), .C(n5460), .D(n5351), .Y(n2332) );
  INVX1 U6560 ( .A(inst_register_registers[110]), .Y(n5330) );
  OAI22X1 U6561 ( .A(n5330), .B(n5345), .C(n5462), .D(n5316), .Y(n2331) );
  INVX1 U6562 ( .A(inst_register_registers[111]), .Y(n5331) );
  OAI22X1 U6563 ( .A(n5331), .B(n5345), .C(n5464), .D(n5316), .Y(n2330) );
  INVX1 U6564 ( .A(inst_register_registers[112]), .Y(n5332) );
  OAI22X1 U6565 ( .A(n5332), .B(n5345), .C(n5466), .D(n5351), .Y(n2329) );
  INVX1 U6566 ( .A(inst_register_registers[113]), .Y(n5333) );
  OAI22X1 U6567 ( .A(n5333), .B(n5345), .C(n5468), .D(n5316), .Y(n2328) );
  INVX1 U6568 ( .A(inst_register_registers[114]), .Y(n5334) );
  OAI22X1 U6569 ( .A(n5334), .B(n5345), .C(n5470), .D(n5316), .Y(n2327) );
  INVX1 U6570 ( .A(inst_register_registers[115]), .Y(n5335) );
  OAI22X1 U6571 ( .A(n5335), .B(n5345), .C(n5472), .D(n5351), .Y(n2326) );
  INVX1 U6572 ( .A(inst_register_registers[116]), .Y(n5336) );
  OAI22X1 U6573 ( .A(n5336), .B(n5345), .C(n5474), .D(n5316), .Y(n2325) );
  INVX1 U6574 ( .A(inst_register_registers[117]), .Y(n5337) );
  OAI22X1 U6575 ( .A(n5337), .B(n5317), .C(n5476), .D(n5351), .Y(n2324) );
  INVX1 U6576 ( .A(inst_register_registers[118]), .Y(n5338) );
  OAI22X1 U6577 ( .A(n5338), .B(n5345), .C(n5478), .D(n5316), .Y(n2323) );
  INVX1 U6578 ( .A(inst_register_registers[119]), .Y(n5339) );
  OAI22X1 U6579 ( .A(n5339), .B(n5345), .C(n5480), .D(n5351), .Y(n2322) );
  INVX1 U6580 ( .A(inst_register_registers[120]), .Y(n5340) );
  OAI22X1 U6581 ( .A(n5340), .B(n5345), .C(n5482), .D(n5351), .Y(n2321) );
  INVX1 U6582 ( .A(inst_register_registers[121]), .Y(n5341) );
  OAI22X1 U6583 ( .A(n5341), .B(n5345), .C(n5484), .D(n5316), .Y(n2320) );
  INVX1 U6584 ( .A(inst_register_registers[122]), .Y(n5342) );
  OAI22X1 U6585 ( .A(n5342), .B(n5317), .C(n5487), .D(n5316), .Y(n2319) );
  INVX1 U6586 ( .A(inst_register_registers[123]), .Y(n5343) );
  OAI22X1 U6587 ( .A(n5343), .B(n5317), .C(n5489), .D(n5316), .Y(n2318) );
  INVX1 U6588 ( .A(inst_register_registers[124]), .Y(n5344) );
  OAI22X1 U6589 ( .A(n5344), .B(n5317), .C(n5491), .D(n5316), .Y(n2317) );
  INVX1 U6590 ( .A(inst_register_registers[125]), .Y(n5346) );
  OAI22X1 U6591 ( .A(n5346), .B(n5345), .C(n5493), .D(n5316), .Y(n2316) );
  INVX1 U6592 ( .A(inst_register_registers[126]), .Y(n5347) );
  OAI22X1 U6593 ( .A(n5347), .B(n5317), .C(n5495), .D(n5351), .Y(n2315) );
  INVX1 U6594 ( .A(inst_register_registers[255]), .Y(n5348) );
  OAI22X1 U6595 ( .A(n5348), .B(n2811), .C(n5120), .D(n5431), .Y(n2314) );
  INVX1 U6596 ( .A(inst_register_registers[98]), .Y(n5349) );
  OAI22X1 U6597 ( .A(n5349), .B(n5317), .C(n5438), .D(n5316), .Y(n2313) );
  INVX1 U6598 ( .A(inst_register_registers[96]), .Y(n5350) );
  OAI22X1 U6599 ( .A(n5350), .B(n5317), .C(n5433), .D(n5351), .Y(n2312) );
  INVX1 U6600 ( .A(inst_register_registers[97]), .Y(n5352) );
  OAI22X1 U6601 ( .A(n5352), .B(n5317), .C(n5435), .D(n5351), .Y(n2311) );
  INVX1 U6602 ( .A(inst_register_registers[95]), .Y(n5356) );
  NOR2X1 U6603 ( .A(reg_write_address_WB[2]), .B(n5353), .Y(n5429) );
  NAND2X1 U6604 ( .A(reg_write_address_WB[1]), .B(n5429), .Y(n5388) );
  NAND2X1 U6605 ( .A(n2815), .B(n5354), .Y(n5386) );
  OAI22X1 U6606 ( .A(n5356), .B(n5355), .C(n5431), .D(n5354), .Y(n2310) );
  INVX1 U6607 ( .A(inst_register_registers[64]), .Y(n5357) );
  OAI22X1 U6608 ( .A(n5357), .B(n5355), .C(n5433), .D(n5354), .Y(n2309) );
  INVX1 U6609 ( .A(inst_register_registers[65]), .Y(n5358) );
  OAI22X1 U6610 ( .A(n5358), .B(n5355), .C(n5435), .D(n5354), .Y(n2308) );
  INVX1 U6611 ( .A(inst_register_registers[66]), .Y(n5359) );
  OAI22X1 U6612 ( .A(n5359), .B(n5355), .C(n5438), .D(n5354), .Y(n2307) );
  INVX1 U6613 ( .A(inst_register_registers[67]), .Y(n5360) );
  OAI22X1 U6614 ( .A(n5360), .B(n5355), .C(n5440), .D(n5354), .Y(n2306) );
  INVX1 U6615 ( .A(inst_register_registers[68]), .Y(n5361) );
  OAI22X1 U6616 ( .A(n5361), .B(n5355), .C(n5442), .D(n5354), .Y(n2305) );
  INVX1 U6617 ( .A(inst_register_registers[69]), .Y(n5362) );
  OAI22X1 U6618 ( .A(n5362), .B(n5355), .C(n5444), .D(n5354), .Y(n2304) );
  INVX1 U6619 ( .A(inst_register_registers[70]), .Y(n5363) );
  OAI22X1 U6620 ( .A(n5363), .B(n5355), .C(n5446), .D(n5354), .Y(n2303) );
  INVX1 U6621 ( .A(inst_register_registers[71]), .Y(n5364) );
  OAI22X1 U6622 ( .A(n5364), .B(n5355), .C(n5448), .D(n5388), .Y(n2302) );
  INVX1 U6623 ( .A(inst_register_registers[72]), .Y(n5365) );
  OAI22X1 U6624 ( .A(n5365), .B(n5355), .C(n5450), .D(n5388), .Y(n2301) );
  INVX1 U6625 ( .A(inst_register_registers[73]), .Y(n5366) );
  OAI22X1 U6626 ( .A(n5366), .B(n5355), .C(n5452), .D(n5388), .Y(n2300) );
  INVX1 U6627 ( .A(inst_register_registers[74]), .Y(n5367) );
  OAI22X1 U6628 ( .A(n5367), .B(n5355), .C(n5454), .D(n5388), .Y(n2299) );
  INVX1 U6629 ( .A(inst_register_registers[75]), .Y(n5368) );
  OAI22X1 U6630 ( .A(n5368), .B(n5386), .C(n5456), .D(n5388), .Y(n2298) );
  INVX1 U6631 ( .A(inst_register_registers[76]), .Y(n5369) );
  OAI22X1 U6632 ( .A(n5369), .B(n5386), .C(n5458), .D(n5388), .Y(n2297) );
  INVX1 U6633 ( .A(inst_register_registers[77]), .Y(n5370) );
  OAI22X1 U6634 ( .A(n5370), .B(n5386), .C(n5460), .D(n5388), .Y(n2296) );
  INVX1 U6635 ( .A(inst_register_registers[78]), .Y(n5371) );
  OAI22X1 U6636 ( .A(n5371), .B(n5386), .C(n5462), .D(n5354), .Y(n2295) );
  INVX1 U6637 ( .A(inst_register_registers[79]), .Y(n5372) );
  OAI22X1 U6638 ( .A(n5372), .B(n5386), .C(n5464), .D(n5354), .Y(n2294) );
  INVX1 U6639 ( .A(inst_register_registers[80]), .Y(n5373) );
  OAI22X1 U6640 ( .A(n5373), .B(n5386), .C(n5466), .D(n5388), .Y(n2293) );
  INVX1 U6641 ( .A(inst_register_registers[81]), .Y(n5374) );
  OAI22X1 U6642 ( .A(n5374), .B(n5386), .C(n5468), .D(n5354), .Y(n2292) );
  INVX1 U6643 ( .A(inst_register_registers[82]), .Y(n5375) );
  OAI22X1 U6644 ( .A(n5375), .B(n5386), .C(n5470), .D(n5354), .Y(n2291) );
  INVX1 U6645 ( .A(inst_register_registers[83]), .Y(n5376) );
  OAI22X1 U6646 ( .A(n5376), .B(n5386), .C(n5472), .D(n5354), .Y(n2290) );
  INVX1 U6647 ( .A(inst_register_registers[84]), .Y(n5377) );
  OAI22X1 U6648 ( .A(n5377), .B(n5386), .C(n5474), .D(n5354), .Y(n2289) );
  INVX1 U6649 ( .A(inst_register_registers[85]), .Y(n5378) );
  OAI22X1 U6650 ( .A(n5378), .B(n5355), .C(n5476), .D(n5354), .Y(n2288) );
  INVX1 U6651 ( .A(inst_register_registers[86]), .Y(n5379) );
  OAI22X1 U6652 ( .A(n5379), .B(n5386), .C(n5478), .D(n5354), .Y(n2287) );
  INVX1 U6653 ( .A(inst_register_registers[87]), .Y(n5380) );
  OAI22X1 U6654 ( .A(n5380), .B(n5355), .C(n5480), .D(n5388), .Y(n2286) );
  INVX1 U6655 ( .A(inst_register_registers[88]), .Y(n5381) );
  OAI22X1 U6656 ( .A(n5381), .B(n5355), .C(n5482), .D(n5388), .Y(n2285) );
  INVX1 U6657 ( .A(inst_register_registers[89]), .Y(n5382) );
  OAI22X1 U6658 ( .A(n5382), .B(n5355), .C(n5484), .D(n5354), .Y(n2284) );
  INVX1 U6659 ( .A(inst_register_registers[90]), .Y(n5383) );
  OAI22X1 U6660 ( .A(n5383), .B(n5355), .C(n5487), .D(n5388), .Y(n2283) );
  INVX1 U6661 ( .A(inst_register_registers[91]), .Y(n5384) );
  OAI22X1 U6662 ( .A(n5384), .B(n5355), .C(n5489), .D(n5354), .Y(n2282) );
  INVX1 U6663 ( .A(inst_register_registers[92]), .Y(n5385) );
  OAI22X1 U6664 ( .A(n5385), .B(n5355), .C(n5491), .D(n5354), .Y(n2281) );
  INVX1 U6665 ( .A(inst_register_registers[93]), .Y(n5387) );
  OAI22X1 U6666 ( .A(n5387), .B(n5386), .C(n5493), .D(n5354), .Y(n2280) );
  INVX1 U6667 ( .A(inst_register_registers[94]), .Y(n5389) );
  OAI22X1 U6668 ( .A(n5389), .B(n5355), .C(n5495), .D(n5388), .Y(n2279) );
  OAI21X1 U6669 ( .A(n5392), .B(n5391), .C(n5390), .Y(n5393) );
  INVX1 U6670 ( .A(inst_register_registers[63]), .Y(n5394) );
  AOI22X1 U6671 ( .A(n5427), .B(n5431), .C(n5394), .D(n5425), .Y(n2278) );
  INVX1 U6672 ( .A(inst_register_registers[32]), .Y(n5395) );
  AOI22X1 U6673 ( .A(n5427), .B(n5433), .C(n5395), .D(n5425), .Y(n2277) );
  INVX1 U6674 ( .A(inst_register_registers[33]), .Y(n5396) );
  AOI22X1 U6675 ( .A(n5427), .B(n5435), .C(n5396), .D(n5425), .Y(n2276) );
  INVX1 U6676 ( .A(inst_register_registers[34]), .Y(n5397) );
  AOI22X1 U6677 ( .A(n5427), .B(n5438), .C(n5397), .D(n5425), .Y(n2275) );
  INVX1 U6678 ( .A(inst_register_registers[35]), .Y(n5398) );
  AOI22X1 U6679 ( .A(n5427), .B(n5440), .C(n5398), .D(n5425), .Y(n2274) );
  INVX1 U6680 ( .A(inst_register_registers[36]), .Y(n5399) );
  AOI22X1 U6681 ( .A(n5427), .B(n5442), .C(n5399), .D(n5425), .Y(n2273) );
  INVX1 U6682 ( .A(inst_register_registers[37]), .Y(n5400) );
  AOI22X1 U6683 ( .A(n5427), .B(n5444), .C(n5400), .D(n5425), .Y(n2272) );
  INVX1 U6684 ( .A(inst_register_registers[38]), .Y(n5401) );
  AOI22X1 U6685 ( .A(n5427), .B(n5446), .C(n5401), .D(n5425), .Y(n2271) );
  INVX1 U6686 ( .A(inst_register_registers[39]), .Y(n5402) );
  AOI22X1 U6687 ( .A(n5427), .B(n5448), .C(n5402), .D(n5425), .Y(n2270) );
  INVX1 U6688 ( .A(inst_register_registers[40]), .Y(n5403) );
  AOI22X1 U6689 ( .A(n5427), .B(n5450), .C(n5403), .D(n5425), .Y(n2269) );
  INVX1 U6690 ( .A(inst_register_registers[41]), .Y(n5404) );
  AOI22X1 U6691 ( .A(n5427), .B(n5452), .C(n5404), .D(n5425), .Y(n2268) );
  INVX1 U6692 ( .A(inst_register_registers[42]), .Y(n5405) );
  AOI22X1 U6693 ( .A(n5427), .B(n5454), .C(n5405), .D(n5425), .Y(n2267) );
  INVX1 U6694 ( .A(inst_register_registers[43]), .Y(n5406) );
  AOI22X1 U6695 ( .A(n5427), .B(n5456), .C(n5406), .D(n5425), .Y(n2266) );
  INVX1 U6696 ( .A(inst_register_registers[44]), .Y(n5407) );
  AOI22X1 U6697 ( .A(n5427), .B(n5458), .C(n5407), .D(n5425), .Y(n2265) );
  INVX1 U6698 ( .A(inst_register_registers[45]), .Y(n5408) );
  AOI22X1 U6699 ( .A(n5427), .B(n5460), .C(n5408), .D(n5425), .Y(n2264) );
  INVX1 U6700 ( .A(inst_register_registers[46]), .Y(n5409) );
  AOI22X1 U6701 ( .A(n5427), .B(n5462), .C(n5409), .D(n5425), .Y(n2263) );
  INVX1 U6702 ( .A(inst_register_registers[47]), .Y(n5410) );
  AOI22X1 U6703 ( .A(n5427), .B(n5464), .C(n5410), .D(n5425), .Y(n2262) );
  INVX1 U6704 ( .A(inst_register_registers[48]), .Y(n5411) );
  AOI22X1 U6705 ( .A(n5427), .B(n5466), .C(n5411), .D(n5425), .Y(n2261) );
  INVX1 U6706 ( .A(inst_register_registers[49]), .Y(n5412) );
  AOI22X1 U6707 ( .A(n5427), .B(n5468), .C(n5412), .D(n5425), .Y(n2260) );
  INVX1 U6708 ( .A(inst_register_registers[50]), .Y(n5413) );
  AOI22X1 U6709 ( .A(n5427), .B(n5470), .C(n5413), .D(n5393), .Y(n2259) );
  INVX1 U6710 ( .A(inst_register_registers[51]), .Y(n5414) );
  AOI22X1 U6711 ( .A(n5427), .B(n5472), .C(n5414), .D(n5393), .Y(n2258) );
  INVX1 U6712 ( .A(inst_register_registers[52]), .Y(n5415) );
  AOI22X1 U6713 ( .A(n5427), .B(n5474), .C(n5415), .D(n5393), .Y(n2257) );
  INVX1 U6714 ( .A(inst_register_registers[53]), .Y(n5416) );
  AOI22X1 U6715 ( .A(n5427), .B(n5476), .C(n5416), .D(n5393), .Y(n2256) );
  INVX1 U6716 ( .A(inst_register_registers[54]), .Y(n5417) );
  AOI22X1 U6717 ( .A(n5427), .B(n5478), .C(n5417), .D(n5425), .Y(n2255) );
  INVX1 U6718 ( .A(inst_register_registers[55]), .Y(n5418) );
  AOI22X1 U6719 ( .A(n5427), .B(n5480), .C(n5418), .D(n5393), .Y(n2254) );
  INVX1 U6720 ( .A(inst_register_registers[56]), .Y(n5419) );
  AOI22X1 U6721 ( .A(n5427), .B(n5482), .C(n5419), .D(n5425), .Y(n2253) );
  INVX1 U6722 ( .A(inst_register_registers[57]), .Y(n5420) );
  INVX2 U6723 ( .A(n5427), .Y(n5425) );
  AOI22X1 U6724 ( .A(n5427), .B(n5484), .C(n5420), .D(n5425), .Y(n2252) );
  INVX1 U6725 ( .A(inst_register_registers[58]), .Y(n5421) );
  AOI22X1 U6726 ( .A(n5427), .B(n5487), .C(n5421), .D(n5425), .Y(n2251) );
  INVX1 U6727 ( .A(inst_register_registers[59]), .Y(n5422) );
  AOI22X1 U6728 ( .A(n5427), .B(n5489), .C(n5422), .D(n5425), .Y(n2250) );
  INVX1 U6729 ( .A(inst_register_registers[60]), .Y(n5423) );
  AOI22X1 U6730 ( .A(n5427), .B(n5491), .C(n5423), .D(n5425), .Y(n2249) );
  INVX1 U6731 ( .A(inst_register_registers[61]), .Y(n5424) );
  AOI22X1 U6732 ( .A(n5427), .B(n5493), .C(n5424), .D(n5425), .Y(n2248) );
  INVX1 U6733 ( .A(inst_register_registers[62]), .Y(n5426) );
  AOI22X1 U6734 ( .A(n5427), .B(n5495), .C(n5426), .D(n5425), .Y(n2247) );
  INVX1 U6735 ( .A(inst_register_registers[31]), .Y(n5432) );
  NAND2X1 U6736 ( .A(n5429), .B(n5428), .Y(n5486) );
  AND2X2 U6737 ( .A(n3066), .B(n5430), .Y(n5437) );
  OAI22X1 U6738 ( .A(n5432), .B(n2813), .C(n5431), .D(n5430), .Y(n2246) );
  INVX1 U6739 ( .A(inst_register_registers[0]), .Y(n5434) );
  OAI22X1 U6740 ( .A(n5434), .B(n2813), .C(n5433), .D(n5430), .Y(n2245) );
  INVX1 U6741 ( .A(inst_register_registers[1]), .Y(n5436) );
  OAI22X1 U6742 ( .A(n5436), .B(n2813), .C(n5435), .D(n5430), .Y(n2244) );
  INVX1 U6743 ( .A(inst_register_registers[2]), .Y(n5439) );
  OAI22X1 U6744 ( .A(n5439), .B(n2813), .C(n5438), .D(n5430), .Y(n2243) );
  INVX1 U6745 ( .A(inst_register_registers[3]), .Y(n5441) );
  OAI22X1 U6746 ( .A(n5441), .B(n2813), .C(n5440), .D(n5430), .Y(n2242) );
  INVX1 U6747 ( .A(inst_register_registers[4]), .Y(n5443) );
  OAI22X1 U6748 ( .A(n5443), .B(n2813), .C(n5442), .D(n5430), .Y(n2241) );
  INVX1 U6749 ( .A(inst_register_registers[5]), .Y(n5445) );
  OAI22X1 U6750 ( .A(n5445), .B(n2813), .C(n5444), .D(n5430), .Y(n2240) );
  INVX1 U6751 ( .A(inst_register_registers[6]), .Y(n5447) );
  OAI22X1 U6752 ( .A(n5447), .B(n2813), .C(n5446), .D(n5486), .Y(n2239) );
  INVX1 U6753 ( .A(inst_register_registers[7]), .Y(n5449) );
  OAI22X1 U6754 ( .A(n5449), .B(n2813), .C(n5448), .D(n5486), .Y(n2238) );
  INVX1 U6755 ( .A(inst_register_registers[8]), .Y(n5451) );
  OAI22X1 U6756 ( .A(n5451), .B(n2813), .C(n5450), .D(n5486), .Y(n2237) );
  INVX1 U6757 ( .A(inst_register_registers[9]), .Y(n5453) );
  OAI22X1 U6758 ( .A(n5453), .B(n2813), .C(n5452), .D(n5486), .Y(n2236) );
  INVX1 U6759 ( .A(inst_register_registers[10]), .Y(n5455) );
  OAI22X1 U6760 ( .A(n5455), .B(n2813), .C(n5454), .D(n5486), .Y(n2235) );
  INVX1 U6761 ( .A(inst_register_registers[11]), .Y(n5457) );
  OAI22X1 U6762 ( .A(n5457), .B(n2813), .C(n5456), .D(n5486), .Y(n2234) );
  INVX1 U6763 ( .A(inst_register_registers[12]), .Y(n5459) );
  OAI22X1 U6764 ( .A(n5459), .B(n2813), .C(n5458), .D(n5430), .Y(n2233) );
  INVX1 U6765 ( .A(inst_register_registers[13]), .Y(n5461) );
  OAI22X1 U6766 ( .A(n5461), .B(n2813), .C(n5460), .D(n5430), .Y(n2232) );
  INVX1 U6767 ( .A(inst_register_registers[14]), .Y(n5463) );
  OAI22X1 U6768 ( .A(n5463), .B(n2813), .C(n5462), .D(n5430), .Y(n2231) );
  INVX1 U6769 ( .A(inst_register_registers[15]), .Y(n5465) );
  OAI22X1 U6770 ( .A(n5465), .B(n2813), .C(n5464), .D(n5430), .Y(n2230) );
  INVX1 U6771 ( .A(inst_register_registers[16]), .Y(n5467) );
  OAI22X1 U6772 ( .A(n5467), .B(n2813), .C(n5466), .D(n5486), .Y(n2229) );
  INVX1 U6773 ( .A(inst_register_registers[17]), .Y(n5469) );
  OAI22X1 U6774 ( .A(n5469), .B(n2813), .C(n5468), .D(n5430), .Y(n2228) );
  INVX1 U6775 ( .A(inst_register_registers[18]), .Y(n5471) );
  OAI22X1 U6776 ( .A(n5471), .B(n2813), .C(n5470), .D(n5430), .Y(n2227) );
  INVX1 U6777 ( .A(inst_register_registers[19]), .Y(n5473) );
  OAI22X1 U6778 ( .A(n5473), .B(n2813), .C(n5472), .D(n5430), .Y(n2226) );
  INVX1 U6779 ( .A(inst_register_registers[20]), .Y(n5475) );
  OAI22X1 U6780 ( .A(n5475), .B(n2813), .C(n5474), .D(n5486), .Y(n2225) );
  INVX1 U6781 ( .A(inst_register_registers[21]), .Y(n5477) );
  OAI22X1 U6782 ( .A(n5477), .B(n2813), .C(n5476), .D(n5430), .Y(n2224) );
  INVX1 U6783 ( .A(inst_register_registers[22]), .Y(n5479) );
  OAI22X1 U6784 ( .A(n5479), .B(n2813), .C(n5478), .D(n5486), .Y(n2223) );
  INVX1 U6785 ( .A(inst_register_registers[23]), .Y(n5481) );
  AOI22X1 U6786 ( .A(n5481), .B(n5430), .C(n5480), .D(n2813), .Y(n2222) );
  INVX1 U6787 ( .A(inst_register_registers[24]), .Y(n5483) );
  OAI22X1 U6788 ( .A(n5483), .B(n2813), .C(n5482), .D(n5486), .Y(n2221) );
  INVX1 U6789 ( .A(inst_register_registers[25]), .Y(n5485) );
  OAI22X1 U6790 ( .A(n5485), .B(n2813), .C(n5484), .D(n5486), .Y(n2220) );
  INVX1 U6791 ( .A(inst_register_registers[26]), .Y(n5488) );
  OAI22X1 U6792 ( .A(n5488), .B(n2813), .C(n5487), .D(n5486), .Y(n2219) );
  INVX1 U6793 ( .A(inst_register_registers[27]), .Y(n5490) );
  OAI22X1 U6794 ( .A(n5490), .B(n2813), .C(n5489), .D(n5430), .Y(n2218) );
  INVX1 U6795 ( .A(inst_register_registers[28]), .Y(n5492) );
  OAI22X1 U6796 ( .A(n5492), .B(n2813), .C(n5491), .D(n5430), .Y(n2217) );
  INVX1 U6797 ( .A(inst_register_registers[29]), .Y(n5494) );
  OAI22X1 U6798 ( .A(n5494), .B(n2813), .C(n5493), .D(n5430), .Y(n2216) );
  INVX1 U6799 ( .A(inst_register_registers[30]), .Y(n5496) );
  OAI22X1 U6800 ( .A(n5496), .B(n2813), .C(n5495), .D(n5430), .Y(n2215) );
  NAND2X1 U6801 ( .A(n5497), .B(jump_inst_addr_MEM[2]), .Y(n5498) );
  OAI21X1 U6802 ( .A(inst_address[2]), .B(n5524), .C(n5498), .Y(n5499) );
  AOI21X1 U6803 ( .A(n5526), .B(shifted_address_MEM[2]), .C(n5499), .Y(n5500)
         );
  OAI21X1 U6804 ( .A(n5502), .B(n5501), .C(n5500), .Y(n2212) );
  NOR2X1 U6805 ( .A(inst_address[26]), .B(n5524), .Y(n5508) );
  OAI21X1 U6806 ( .A(inst_address[25]), .B(n5524), .C(n5503), .Y(n5507) );
  AOI22X1 U6807 ( .A(inst_address[26]), .B(n5507), .C(n5526), .D(
        shifted_address_MEM[26]), .Y(n5504) );
  OAI21X1 U6808 ( .A(n5506), .B(n5505), .C(n5504), .Y(n2188) );
  NOR2X1 U6809 ( .A(n5508), .B(n5507), .Y(n5513) );
  NOR2X1 U6810 ( .A(inst_address[27]), .B(n5524), .Y(n5510) );
  AOI22X1 U6811 ( .A(n5510), .B(n5509), .C(n5526), .D(shifted_address_MEM[27]), 
        .Y(n5511) );
  OAI21X1 U6812 ( .A(n5513), .B(n5512), .C(n5511), .Y(n2187) );
  NOR2X1 U6813 ( .A(inst_address[28]), .B(n5524), .Y(n5518) );
  OAI21X1 U6814 ( .A(inst_address[27]), .B(n5524), .C(n5513), .Y(n5517) );
  AOI22X1 U6815 ( .A(inst_address[28]), .B(n5517), .C(n5526), .D(
        shifted_address_MEM[28]), .Y(n5514) );
  OAI21X1 U6816 ( .A(n5516), .B(n5515), .C(n5514), .Y(n2186) );
  NOR2X1 U6817 ( .A(n5518), .B(n5517), .Y(n5523) );
  NOR2X1 U6818 ( .A(inst_address[29]), .B(n5524), .Y(n5520) );
  AOI22X1 U6819 ( .A(n5520), .B(n5519), .C(n5526), .D(shifted_address_MEM[29]), 
        .Y(n5521) );
  OAI21X1 U6820 ( .A(n5523), .B(n5522), .C(n5521), .Y(n2185) );
  OAI21X1 U6821 ( .A(inst_address[29]), .B(n5524), .C(n5523), .Y(n5525) );
  AOI22X1 U6822 ( .A(shifted_address_MEM[30]), .B(n5526), .C(inst_address[30]), 
        .D(n5525), .Y(n5527) );
  OAI21X1 U6823 ( .A(inst_address[30]), .B(n5528), .C(n5527), .Y(n2183) );
endmodule
